
module register_file_DATA_WIDTH64_LOG2_NUM_REGS5_NUM_REGS32 ( clk, reset_n, 
        read_en, write_en, raddr_0, raddr_1, waddr, wdata, rdata_0, rdata_1 );
  input [1:0] read_en;
  input [4:0] raddr_0;
  input [4:0] raddr_1;
  input [4:0] waddr;
  input [63:0] wdata;
  output [63:0] rdata_0;
  output [63:0] rdata_1;
  input clk, reset_n, write_en;
  wire   N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, \RF[0][63] ,
         \RF[0][62] , \RF[0][61] , \RF[0][60] , \RF[0][59] , \RF[0][58] ,
         \RF[0][57] , \RF[0][56] , \RF[0][55] , \RF[0][54] , \RF[0][53] ,
         \RF[0][52] , \RF[0][51] , \RF[0][50] , \RF[0][49] , \RF[0][48] ,
         \RF[0][47] , \RF[0][46] , \RF[0][45] , \RF[0][44] , \RF[0][43] ,
         \RF[0][42] , \RF[0][41] , \RF[0][40] , \RF[0][39] , \RF[0][38] ,
         \RF[0][37] , \RF[0][36] , \RF[0][35] , \RF[0][34] , \RF[0][33] ,
         \RF[0][32] , \RF[0][31] , \RF[0][30] , \RF[0][29] , \RF[0][28] ,
         \RF[0][27] , \RF[0][26] , \RF[0][25] , \RF[0][24] , \RF[0][23] ,
         \RF[0][22] , \RF[0][21] , \RF[0][20] , \RF[0][19] , \RF[0][18] ,
         \RF[0][17] , \RF[0][16] , \RF[0][15] , \RF[0][14] , \RF[0][13] ,
         \RF[0][12] , \RF[0][11] , \RF[0][10] , \RF[0][9] , \RF[0][8] ,
         \RF[0][7] , \RF[0][6] , \RF[0][5] , \RF[0][4] , \RF[0][3] ,
         \RF[0][2] , \RF[0][1] , \RF[0][0] , \RF[1][63] , \RF[1][62] ,
         \RF[1][61] , \RF[1][60] , \RF[1][59] , \RF[1][58] , \RF[1][57] ,
         \RF[1][56] , \RF[1][55] , \RF[1][54] , \RF[1][53] , \RF[1][52] ,
         \RF[1][51] , \RF[1][50] , \RF[1][49] , \RF[1][48] , \RF[1][47] ,
         \RF[1][46] , \RF[1][45] , \RF[1][44] , \RF[1][43] , \RF[1][42] ,
         \RF[1][41] , \RF[1][40] , \RF[1][39] , \RF[1][38] , \RF[1][37] ,
         \RF[1][36] , \RF[1][35] , \RF[1][34] , \RF[1][33] , \RF[1][32] ,
         \RF[1][31] , \RF[1][30] , \RF[1][29] , \RF[1][28] , \RF[1][27] ,
         \RF[1][26] , \RF[1][25] , \RF[1][24] , \RF[1][23] , \RF[1][22] ,
         \RF[1][21] , \RF[1][20] , \RF[1][19] , \RF[1][18] , \RF[1][17] ,
         \RF[1][16] , \RF[1][15] , \RF[1][14] , \RF[1][13] , \RF[1][12] ,
         \RF[1][11] , \RF[1][10] , \RF[1][9] , \RF[1][8] , \RF[1][7] ,
         \RF[1][6] , \RF[1][5] , \RF[1][4] , \RF[1][3] , \RF[1][2] ,
         \RF[1][1] , \RF[1][0] , \RF[2][63] , \RF[2][62] , \RF[2][61] ,
         \RF[2][60] , \RF[2][59] , \RF[2][58] , \RF[2][57] , \RF[2][56] ,
         \RF[2][55] , \RF[2][54] , \RF[2][53] , \RF[2][52] , \RF[2][51] ,
         \RF[2][50] , \RF[2][49] , \RF[2][48] , \RF[2][47] , \RF[2][46] ,
         \RF[2][45] , \RF[2][44] , \RF[2][43] , \RF[2][42] , \RF[2][41] ,
         \RF[2][40] , \RF[2][39] , \RF[2][38] , \RF[2][37] , \RF[2][36] ,
         \RF[2][35] , \RF[2][34] , \RF[2][33] , \RF[2][32] , \RF[2][31] ,
         \RF[2][30] , \RF[2][29] , \RF[2][28] , \RF[2][27] , \RF[2][26] ,
         \RF[2][25] , \RF[2][24] , \RF[2][23] , \RF[2][22] , \RF[2][21] ,
         \RF[2][20] , \RF[2][19] , \RF[2][18] , \RF[2][17] , \RF[2][16] ,
         \RF[2][15] , \RF[2][14] , \RF[2][13] , \RF[2][12] , \RF[2][11] ,
         \RF[2][10] , \RF[2][9] , \RF[2][8] , \RF[2][7] , \RF[2][6] ,
         \RF[2][5] , \RF[2][4] , \RF[2][3] , \RF[2][2] , \RF[2][1] ,
         \RF[2][0] , \RF[3][63] , \RF[3][62] , \RF[3][61] , \RF[3][60] ,
         \RF[3][59] , \RF[3][58] , \RF[3][57] , \RF[3][56] , \RF[3][55] ,
         \RF[3][54] , \RF[3][53] , \RF[3][52] , \RF[3][51] , \RF[3][50] ,
         \RF[3][49] , \RF[3][48] , \RF[3][47] , \RF[3][46] , \RF[3][45] ,
         \RF[3][44] , \RF[3][43] , \RF[3][42] , \RF[3][41] , \RF[3][40] ,
         \RF[3][39] , \RF[3][38] , \RF[3][37] , \RF[3][36] , \RF[3][35] ,
         \RF[3][34] , \RF[3][33] , \RF[3][32] , \RF[3][31] , \RF[3][30] ,
         \RF[3][29] , \RF[3][28] , \RF[3][27] , \RF[3][26] , \RF[3][25] ,
         \RF[3][24] , \RF[3][23] , \RF[3][22] , \RF[3][21] , \RF[3][20] ,
         \RF[3][19] , \RF[3][18] , \RF[3][17] , \RF[3][16] , \RF[3][15] ,
         \RF[3][14] , \RF[3][13] , \RF[3][12] , \RF[3][11] , \RF[3][10] ,
         \RF[3][9] , \RF[3][8] , \RF[3][7] , \RF[3][6] , \RF[3][5] ,
         \RF[3][4] , \RF[3][3] , \RF[3][2] , \RF[3][1] , \RF[3][0] ,
         \RF[4][63] , \RF[4][62] , \RF[4][61] , \RF[4][60] , \RF[4][59] ,
         \RF[4][58] , \RF[4][57] , \RF[4][56] , \RF[4][55] , \RF[4][54] ,
         \RF[4][53] , \RF[4][52] , \RF[4][51] , \RF[4][50] , \RF[4][49] ,
         \RF[4][48] , \RF[4][47] , \RF[4][46] , \RF[4][45] , \RF[4][44] ,
         \RF[4][43] , \RF[4][42] , \RF[4][41] , \RF[4][40] , \RF[4][39] ,
         \RF[4][38] , \RF[4][37] , \RF[4][36] , \RF[4][35] , \RF[4][34] ,
         \RF[4][33] , \RF[4][32] , \RF[4][31] , \RF[4][30] , \RF[4][29] ,
         \RF[4][28] , \RF[4][27] , \RF[4][26] , \RF[4][25] , \RF[4][24] ,
         \RF[4][23] , \RF[4][22] , \RF[4][21] , \RF[4][20] , \RF[4][19] ,
         \RF[4][18] , \RF[4][17] , \RF[4][16] , \RF[4][15] , \RF[4][14] ,
         \RF[4][13] , \RF[4][12] , \RF[4][11] , \RF[4][10] , \RF[4][9] ,
         \RF[4][8] , \RF[4][7] , \RF[4][6] , \RF[4][5] , \RF[4][4] ,
         \RF[4][3] , \RF[4][2] , \RF[4][1] , \RF[4][0] , \RF[5][63] ,
         \RF[5][62] , \RF[5][61] , \RF[5][60] , \RF[5][59] , \RF[5][58] ,
         \RF[5][57] , \RF[5][56] , \RF[5][55] , \RF[5][54] , \RF[5][53] ,
         \RF[5][52] , \RF[5][51] , \RF[5][50] , \RF[5][49] , \RF[5][48] ,
         \RF[5][47] , \RF[5][46] , \RF[5][45] , \RF[5][44] , \RF[5][43] ,
         \RF[5][42] , \RF[5][41] , \RF[5][40] , \RF[5][39] , \RF[5][38] ,
         \RF[5][37] , \RF[5][36] , \RF[5][35] , \RF[5][34] , \RF[5][33] ,
         \RF[5][32] , \RF[5][31] , \RF[5][30] , \RF[5][29] , \RF[5][28] ,
         \RF[5][27] , \RF[5][26] , \RF[5][25] , \RF[5][24] , \RF[5][23] ,
         \RF[5][22] , \RF[5][21] , \RF[5][20] , \RF[5][19] , \RF[5][18] ,
         \RF[5][17] , \RF[5][16] , \RF[5][15] , \RF[5][14] , \RF[5][13] ,
         \RF[5][12] , \RF[5][11] , \RF[5][10] , \RF[5][9] , \RF[5][8] ,
         \RF[5][7] , \RF[5][6] , \RF[5][5] , \RF[5][4] , \RF[5][3] ,
         \RF[5][2] , \RF[5][1] , \RF[5][0] , \RF[6][63] , \RF[6][62] ,
         \RF[6][61] , \RF[6][60] , \RF[6][59] , \RF[6][58] , \RF[6][57] ,
         \RF[6][56] , \RF[6][55] , \RF[6][54] , \RF[6][53] , \RF[6][52] ,
         \RF[6][51] , \RF[6][50] , \RF[6][49] , \RF[6][48] , \RF[6][47] ,
         \RF[6][46] , \RF[6][45] , \RF[6][44] , \RF[6][43] , \RF[6][42] ,
         \RF[6][41] , \RF[6][40] , \RF[6][39] , \RF[6][38] , \RF[6][37] ,
         \RF[6][36] , \RF[6][35] , \RF[6][34] , \RF[6][33] , \RF[6][32] ,
         \RF[6][31] , \RF[6][30] , \RF[6][29] , \RF[6][28] , \RF[6][27] ,
         \RF[6][26] , \RF[6][25] , \RF[6][24] , \RF[6][23] , \RF[6][22] ,
         \RF[6][21] , \RF[6][20] , \RF[6][19] , \RF[6][18] , \RF[6][17] ,
         \RF[6][16] , \RF[6][15] , \RF[6][14] , \RF[6][13] , \RF[6][12] ,
         \RF[6][11] , \RF[6][10] , \RF[6][9] , \RF[6][8] , \RF[6][7] ,
         \RF[6][6] , \RF[6][5] , \RF[6][4] , \RF[6][3] , \RF[6][2] ,
         \RF[6][1] , \RF[6][0] , \RF[7][63] , \RF[7][62] , \RF[7][61] ,
         \RF[7][60] , \RF[7][59] , \RF[7][58] , \RF[7][57] , \RF[7][56] ,
         \RF[7][55] , \RF[7][54] , \RF[7][53] , \RF[7][52] , \RF[7][51] ,
         \RF[7][50] , \RF[7][49] , \RF[7][48] , \RF[7][47] , \RF[7][46] ,
         \RF[7][45] , \RF[7][44] , \RF[7][43] , \RF[7][42] , \RF[7][41] ,
         \RF[7][40] , \RF[7][39] , \RF[7][38] , \RF[7][37] , \RF[7][36] ,
         \RF[7][35] , \RF[7][34] , \RF[7][33] , \RF[7][32] , \RF[7][31] ,
         \RF[7][30] , \RF[7][29] , \RF[7][28] , \RF[7][27] , \RF[7][26] ,
         \RF[7][25] , \RF[7][24] , \RF[7][23] , \RF[7][22] , \RF[7][21] ,
         \RF[7][20] , \RF[7][19] , \RF[7][18] , \RF[7][17] , \RF[7][16] ,
         \RF[7][15] , \RF[7][14] , \RF[7][13] , \RF[7][12] , \RF[7][11] ,
         \RF[7][10] , \RF[7][9] , \RF[7][8] , \RF[7][7] , \RF[7][6] ,
         \RF[7][5] , \RF[7][4] , \RF[7][3] , \RF[7][2] , \RF[7][1] ,
         \RF[7][0] , \RF[8][63] , \RF[8][62] , \RF[8][61] , \RF[8][60] ,
         \RF[8][59] , \RF[8][58] , \RF[8][57] , \RF[8][56] , \RF[8][55] ,
         \RF[8][54] , \RF[8][53] , \RF[8][52] , \RF[8][51] , \RF[8][50] ,
         \RF[8][49] , \RF[8][48] , \RF[8][47] , \RF[8][46] , \RF[8][45] ,
         \RF[8][44] , \RF[8][43] , \RF[8][42] , \RF[8][41] , \RF[8][40] ,
         \RF[8][39] , \RF[8][38] , \RF[8][37] , \RF[8][36] , \RF[8][35] ,
         \RF[8][34] , \RF[8][33] , \RF[8][32] , \RF[8][31] , \RF[8][30] ,
         \RF[8][29] , \RF[8][28] , \RF[8][27] , \RF[8][26] , \RF[8][25] ,
         \RF[8][24] , \RF[8][23] , \RF[8][22] , \RF[8][21] , \RF[8][20] ,
         \RF[8][19] , \RF[8][18] , \RF[8][17] , \RF[8][16] , \RF[8][15] ,
         \RF[8][14] , \RF[8][13] , \RF[8][12] , \RF[8][11] , \RF[8][10] ,
         \RF[8][9] , \RF[8][8] , \RF[8][7] , \RF[8][6] , \RF[8][5] ,
         \RF[8][4] , \RF[8][3] , \RF[8][2] , \RF[8][1] , \RF[8][0] ,
         \RF[9][63] , \RF[9][62] , \RF[9][61] , \RF[9][60] , \RF[9][59] ,
         \RF[9][58] , \RF[9][57] , \RF[9][56] , \RF[9][55] , \RF[9][54] ,
         \RF[9][53] , \RF[9][52] , \RF[9][51] , \RF[9][50] , \RF[9][49] ,
         \RF[9][48] , \RF[9][47] , \RF[9][46] , \RF[9][45] , \RF[9][44] ,
         \RF[9][43] , \RF[9][42] , \RF[9][41] , \RF[9][40] , \RF[9][39] ,
         \RF[9][38] , \RF[9][37] , \RF[9][36] , \RF[9][35] , \RF[9][34] ,
         \RF[9][33] , \RF[9][32] , \RF[9][31] , \RF[9][30] , \RF[9][29] ,
         \RF[9][28] , \RF[9][27] , \RF[9][26] , \RF[9][25] , \RF[9][24] ,
         \RF[9][23] , \RF[9][22] , \RF[9][21] , \RF[9][20] , \RF[9][19] ,
         \RF[9][18] , \RF[9][17] , \RF[9][16] , \RF[9][15] , \RF[9][14] ,
         \RF[9][13] , \RF[9][12] , \RF[9][11] , \RF[9][10] , \RF[9][9] ,
         \RF[9][8] , \RF[9][7] , \RF[9][6] , \RF[9][5] , \RF[9][4] ,
         \RF[9][3] , \RF[9][2] , \RF[9][1] , \RF[9][0] , \RF[10][63] ,
         \RF[10][62] , \RF[10][61] , \RF[10][60] , \RF[10][59] , \RF[10][58] ,
         \RF[10][57] , \RF[10][56] , \RF[10][55] , \RF[10][54] , \RF[10][53] ,
         \RF[10][52] , \RF[10][51] , \RF[10][50] , \RF[10][49] , \RF[10][48] ,
         \RF[10][47] , \RF[10][46] , \RF[10][45] , \RF[10][44] , \RF[10][43] ,
         \RF[10][42] , \RF[10][41] , \RF[10][40] , \RF[10][39] , \RF[10][38] ,
         \RF[10][37] , \RF[10][36] , \RF[10][35] , \RF[10][34] , \RF[10][33] ,
         \RF[10][32] , \RF[10][31] , \RF[10][30] , \RF[10][29] , \RF[10][28] ,
         \RF[10][27] , \RF[10][26] , \RF[10][25] , \RF[10][24] , \RF[10][23] ,
         \RF[10][22] , \RF[10][21] , \RF[10][20] , \RF[10][19] , \RF[10][18] ,
         \RF[10][17] , \RF[10][16] , \RF[10][15] , \RF[10][14] , \RF[10][13] ,
         \RF[10][12] , \RF[10][11] , \RF[10][10] , \RF[10][9] , \RF[10][8] ,
         \RF[10][7] , \RF[10][6] , \RF[10][5] , \RF[10][4] , \RF[10][3] ,
         \RF[10][2] , \RF[10][1] , \RF[10][0] , \RF[11][63] , \RF[11][62] ,
         \RF[11][61] , \RF[11][60] , \RF[11][59] , \RF[11][58] , \RF[11][57] ,
         \RF[11][56] , \RF[11][55] , \RF[11][54] , \RF[11][53] , \RF[11][52] ,
         \RF[11][51] , \RF[11][50] , \RF[11][49] , \RF[11][48] , \RF[11][47] ,
         \RF[11][46] , \RF[11][45] , \RF[11][44] , \RF[11][43] , \RF[11][42] ,
         \RF[11][41] , \RF[11][40] , \RF[11][39] , \RF[11][38] , \RF[11][37] ,
         \RF[11][36] , \RF[11][35] , \RF[11][34] , \RF[11][33] , \RF[11][32] ,
         \RF[11][31] , \RF[11][30] , \RF[11][29] , \RF[11][28] , \RF[11][27] ,
         \RF[11][26] , \RF[11][25] , \RF[11][24] , \RF[11][23] , \RF[11][22] ,
         \RF[11][21] , \RF[11][20] , \RF[11][19] , \RF[11][18] , \RF[11][17] ,
         \RF[11][16] , \RF[11][15] , \RF[11][14] , \RF[11][13] , \RF[11][12] ,
         \RF[11][11] , \RF[11][10] , \RF[11][9] , \RF[11][8] , \RF[11][7] ,
         \RF[11][6] , \RF[11][5] , \RF[11][4] , \RF[11][3] , \RF[11][2] ,
         \RF[11][1] , \RF[11][0] , \RF[12][63] , \RF[12][62] , \RF[12][61] ,
         \RF[12][60] , \RF[12][59] , \RF[12][58] , \RF[12][57] , \RF[12][56] ,
         \RF[12][55] , \RF[12][54] , \RF[12][53] , \RF[12][52] , \RF[12][51] ,
         \RF[12][50] , \RF[12][49] , \RF[12][48] , \RF[12][47] , \RF[12][46] ,
         \RF[12][45] , \RF[12][44] , \RF[12][43] , \RF[12][42] , \RF[12][41] ,
         \RF[12][40] , \RF[12][39] , \RF[12][38] , \RF[12][37] , \RF[12][36] ,
         \RF[12][35] , \RF[12][34] , \RF[12][33] , \RF[12][32] , \RF[12][31] ,
         \RF[12][30] , \RF[12][29] , \RF[12][28] , \RF[12][27] , \RF[12][26] ,
         \RF[12][25] , \RF[12][24] , \RF[12][23] , \RF[12][22] , \RF[12][21] ,
         \RF[12][20] , \RF[12][19] , \RF[12][18] , \RF[12][17] , \RF[12][16] ,
         \RF[12][15] , \RF[12][14] , \RF[12][13] , \RF[12][12] , \RF[12][11] ,
         \RF[12][10] , \RF[12][9] , \RF[12][8] , \RF[12][7] , \RF[12][6] ,
         \RF[12][5] , \RF[12][4] , \RF[12][3] , \RF[12][2] , \RF[12][1] ,
         \RF[12][0] , \RF[13][63] , \RF[13][62] , \RF[13][61] , \RF[13][60] ,
         \RF[13][59] , \RF[13][58] , \RF[13][57] , \RF[13][56] , \RF[13][55] ,
         \RF[13][54] , \RF[13][53] , \RF[13][52] , \RF[13][51] , \RF[13][50] ,
         \RF[13][49] , \RF[13][48] , \RF[13][47] , \RF[13][46] , \RF[13][45] ,
         \RF[13][44] , \RF[13][43] , \RF[13][42] , \RF[13][41] , \RF[13][40] ,
         \RF[13][39] , \RF[13][38] , \RF[13][37] , \RF[13][36] , \RF[13][35] ,
         \RF[13][34] , \RF[13][33] , \RF[13][32] , \RF[13][31] , \RF[13][30] ,
         \RF[13][29] , \RF[13][28] , \RF[13][27] , \RF[13][26] , \RF[13][25] ,
         \RF[13][24] , \RF[13][23] , \RF[13][22] , \RF[13][21] , \RF[13][20] ,
         \RF[13][19] , \RF[13][18] , \RF[13][17] , \RF[13][16] , \RF[13][15] ,
         \RF[13][14] , \RF[13][13] , \RF[13][12] , \RF[13][11] , \RF[13][10] ,
         \RF[13][9] , \RF[13][8] , \RF[13][7] , \RF[13][6] , \RF[13][5] ,
         \RF[13][4] , \RF[13][3] , \RF[13][2] , \RF[13][1] , \RF[13][0] ,
         \RF[14][63] , \RF[14][62] , \RF[14][61] , \RF[14][60] , \RF[14][59] ,
         \RF[14][58] , \RF[14][57] , \RF[14][56] , \RF[14][55] , \RF[14][54] ,
         \RF[14][53] , \RF[14][52] , \RF[14][51] , \RF[14][50] , \RF[14][49] ,
         \RF[14][48] , \RF[14][47] , \RF[14][46] , \RF[14][45] , \RF[14][44] ,
         \RF[14][43] , \RF[14][42] , \RF[14][41] , \RF[14][40] , \RF[14][39] ,
         \RF[14][38] , \RF[14][37] , \RF[14][36] , \RF[14][35] , \RF[14][34] ,
         \RF[14][33] , \RF[14][32] , \RF[14][31] , \RF[14][30] , \RF[14][29] ,
         \RF[14][28] , \RF[14][27] , \RF[14][26] , \RF[14][25] , \RF[14][24] ,
         \RF[14][23] , \RF[14][22] , \RF[14][21] , \RF[14][20] , \RF[14][19] ,
         \RF[14][18] , \RF[14][17] , \RF[14][16] , \RF[14][15] , \RF[14][14] ,
         \RF[14][13] , \RF[14][12] , \RF[14][11] , \RF[14][10] , \RF[14][9] ,
         \RF[14][8] , \RF[14][7] , \RF[14][6] , \RF[14][5] , \RF[14][4] ,
         \RF[14][3] , \RF[14][2] , \RF[14][1] , \RF[14][0] , \RF[15][63] ,
         \RF[15][62] , \RF[15][61] , \RF[15][60] , \RF[15][59] , \RF[15][58] ,
         \RF[15][57] , \RF[15][56] , \RF[15][55] , \RF[15][54] , \RF[15][53] ,
         \RF[15][52] , \RF[15][51] , \RF[15][50] , \RF[15][49] , \RF[15][48] ,
         \RF[15][47] , \RF[15][46] , \RF[15][45] , \RF[15][44] , \RF[15][43] ,
         \RF[15][42] , \RF[15][41] , \RF[15][40] , \RF[15][39] , \RF[15][38] ,
         \RF[15][37] , \RF[15][36] , \RF[15][35] , \RF[15][34] , \RF[15][33] ,
         \RF[15][32] , \RF[15][31] , \RF[15][30] , \RF[15][29] , \RF[15][28] ,
         \RF[15][27] , \RF[15][26] , \RF[15][25] , \RF[15][24] , \RF[15][23] ,
         \RF[15][22] , \RF[15][21] , \RF[15][20] , \RF[15][19] , \RF[15][18] ,
         \RF[15][17] , \RF[15][16] , \RF[15][15] , \RF[15][14] , \RF[15][13] ,
         \RF[15][12] , \RF[15][11] , \RF[15][10] , \RF[15][9] , \RF[15][8] ,
         \RF[15][7] , \RF[15][6] , \RF[15][5] , \RF[15][4] , \RF[15][3] ,
         \RF[15][2] , \RF[15][1] , \RF[15][0] , \RF[16][63] , \RF[16][62] ,
         \RF[16][61] , \RF[16][60] , \RF[16][59] , \RF[16][58] , \RF[16][57] ,
         \RF[16][56] , \RF[16][55] , \RF[16][54] , \RF[16][53] , \RF[16][52] ,
         \RF[16][51] , \RF[16][50] , \RF[16][49] , \RF[16][48] , \RF[16][47] ,
         \RF[16][46] , \RF[16][45] , \RF[16][44] , \RF[16][43] , \RF[16][42] ,
         \RF[16][41] , \RF[16][40] , \RF[16][39] , \RF[16][38] , \RF[16][37] ,
         \RF[16][36] , \RF[16][35] , \RF[16][34] , \RF[16][33] , \RF[16][32] ,
         \RF[16][31] , \RF[16][30] , \RF[16][29] , \RF[16][28] , \RF[16][27] ,
         \RF[16][26] , \RF[16][25] , \RF[16][24] , \RF[16][23] , \RF[16][22] ,
         \RF[16][21] , \RF[16][20] , \RF[16][19] , \RF[16][18] , \RF[16][17] ,
         \RF[16][16] , \RF[16][15] , \RF[16][14] , \RF[16][13] , \RF[16][12] ,
         \RF[16][11] , \RF[16][10] , \RF[16][9] , \RF[16][8] , \RF[16][7] ,
         \RF[16][6] , \RF[16][5] , \RF[16][4] , \RF[16][3] , \RF[16][2] ,
         \RF[16][1] , \RF[16][0] , \RF[17][63] , \RF[17][62] , \RF[17][61] ,
         \RF[17][60] , \RF[17][59] , \RF[17][58] , \RF[17][57] , \RF[17][56] ,
         \RF[17][55] , \RF[17][54] , \RF[17][53] , \RF[17][52] , \RF[17][51] ,
         \RF[17][50] , \RF[17][49] , \RF[17][48] , \RF[17][47] , \RF[17][46] ,
         \RF[17][45] , \RF[17][44] , \RF[17][43] , \RF[17][42] , \RF[17][41] ,
         \RF[17][40] , \RF[17][39] , \RF[17][38] , \RF[17][37] , \RF[17][36] ,
         \RF[17][35] , \RF[17][34] , \RF[17][33] , \RF[17][32] , \RF[17][31] ,
         \RF[17][30] , \RF[17][29] , \RF[17][28] , \RF[17][27] , \RF[17][26] ,
         \RF[17][25] , \RF[17][24] , \RF[17][23] , \RF[17][22] , \RF[17][21] ,
         \RF[17][20] , \RF[17][19] , \RF[17][18] , \RF[17][17] , \RF[17][16] ,
         \RF[17][15] , \RF[17][14] , \RF[17][13] , \RF[17][12] , \RF[17][11] ,
         \RF[17][10] , \RF[17][9] , \RF[17][8] , \RF[17][7] , \RF[17][6] ,
         \RF[17][5] , \RF[17][4] , \RF[17][3] , \RF[17][2] , \RF[17][1] ,
         \RF[17][0] , \RF[18][63] , \RF[18][62] , \RF[18][61] , \RF[18][60] ,
         \RF[18][59] , \RF[18][58] , \RF[18][57] , \RF[18][56] , \RF[18][55] ,
         \RF[18][54] , \RF[18][53] , \RF[18][52] , \RF[18][51] , \RF[18][50] ,
         \RF[18][49] , \RF[18][48] , \RF[18][47] , \RF[18][46] , \RF[18][45] ,
         \RF[18][44] , \RF[18][43] , \RF[18][42] , \RF[18][41] , \RF[18][40] ,
         \RF[18][39] , \RF[18][38] , \RF[18][37] , \RF[18][36] , \RF[18][35] ,
         \RF[18][34] , \RF[18][33] , \RF[18][32] , \RF[18][31] , \RF[18][30] ,
         \RF[18][29] , \RF[18][28] , \RF[18][27] , \RF[18][26] , \RF[18][25] ,
         \RF[18][24] , \RF[18][23] , \RF[18][22] , \RF[18][21] , \RF[18][20] ,
         \RF[18][19] , \RF[18][18] , \RF[18][17] , \RF[18][16] , \RF[18][15] ,
         \RF[18][14] , \RF[18][13] , \RF[18][12] , \RF[18][11] , \RF[18][10] ,
         \RF[18][9] , \RF[18][8] , \RF[18][7] , \RF[18][6] , \RF[18][5] ,
         \RF[18][4] , \RF[18][3] , \RF[18][2] , \RF[18][1] , \RF[18][0] ,
         \RF[19][63] , \RF[19][62] , \RF[19][61] , \RF[19][60] , \RF[19][59] ,
         \RF[19][58] , \RF[19][57] , \RF[19][56] , \RF[19][55] , \RF[19][54] ,
         \RF[19][53] , \RF[19][52] , \RF[19][51] , \RF[19][50] , \RF[19][49] ,
         \RF[19][48] , \RF[19][47] , \RF[19][46] , \RF[19][45] , \RF[19][44] ,
         \RF[19][43] , \RF[19][42] , \RF[19][41] , \RF[19][40] , \RF[19][39] ,
         \RF[19][38] , \RF[19][37] , \RF[19][36] , \RF[19][35] , \RF[19][34] ,
         \RF[19][33] , \RF[19][32] , \RF[19][31] , \RF[19][30] , \RF[19][29] ,
         \RF[19][28] , \RF[19][27] , \RF[19][26] , \RF[19][25] , \RF[19][24] ,
         \RF[19][23] , \RF[19][22] , \RF[19][21] , \RF[19][20] , \RF[19][19] ,
         \RF[19][18] , \RF[19][17] , \RF[19][16] , \RF[19][15] , \RF[19][14] ,
         \RF[19][13] , \RF[19][12] , \RF[19][11] , \RF[19][10] , \RF[19][9] ,
         \RF[19][8] , \RF[19][7] , \RF[19][6] , \RF[19][5] , \RF[19][4] ,
         \RF[19][3] , \RF[19][2] , \RF[19][1] , \RF[19][0] , \RF[20][63] ,
         \RF[20][62] , \RF[20][61] , \RF[20][60] , \RF[20][59] , \RF[20][58] ,
         \RF[20][57] , \RF[20][56] , \RF[20][55] , \RF[20][54] , \RF[20][53] ,
         \RF[20][52] , \RF[20][51] , \RF[20][50] , \RF[20][49] , \RF[20][48] ,
         \RF[20][47] , \RF[20][46] , \RF[20][45] , \RF[20][44] , \RF[20][43] ,
         \RF[20][42] , \RF[20][41] , \RF[20][40] , \RF[20][39] , \RF[20][38] ,
         \RF[20][37] , \RF[20][36] , \RF[20][35] , \RF[20][34] , \RF[20][33] ,
         \RF[20][32] , \RF[20][31] , \RF[20][30] , \RF[20][29] , \RF[20][28] ,
         \RF[20][27] , \RF[20][26] , \RF[20][25] , \RF[20][24] , \RF[20][23] ,
         \RF[20][22] , \RF[20][21] , \RF[20][20] , \RF[20][19] , \RF[20][18] ,
         \RF[20][17] , \RF[20][16] , \RF[20][15] , \RF[20][14] , \RF[20][13] ,
         \RF[20][12] , \RF[20][11] , \RF[20][10] , \RF[20][9] , \RF[20][8] ,
         \RF[20][7] , \RF[20][6] , \RF[20][5] , \RF[20][4] , \RF[20][3] ,
         \RF[20][2] , \RF[20][1] , \RF[20][0] , \RF[21][63] , \RF[21][62] ,
         \RF[21][61] , \RF[21][60] , \RF[21][59] , \RF[21][58] , \RF[21][57] ,
         \RF[21][56] , \RF[21][55] , \RF[21][54] , \RF[21][53] , \RF[21][52] ,
         \RF[21][51] , \RF[21][50] , \RF[21][49] , \RF[21][48] , \RF[21][47] ,
         \RF[21][46] , \RF[21][45] , \RF[21][44] , \RF[21][43] , \RF[21][42] ,
         \RF[21][41] , \RF[21][40] , \RF[21][39] , \RF[21][38] , \RF[21][37] ,
         \RF[21][36] , \RF[21][35] , \RF[21][34] , \RF[21][33] , \RF[21][32] ,
         \RF[21][31] , \RF[21][30] , \RF[21][29] , \RF[21][28] , \RF[21][27] ,
         \RF[21][26] , \RF[21][25] , \RF[21][24] , \RF[21][23] , \RF[21][22] ,
         \RF[21][21] , \RF[21][20] , \RF[21][19] , \RF[21][18] , \RF[21][17] ,
         \RF[21][16] , \RF[21][15] , \RF[21][14] , \RF[21][13] , \RF[21][12] ,
         \RF[21][11] , \RF[21][10] , \RF[21][9] , \RF[21][8] , \RF[21][7] ,
         \RF[21][6] , \RF[21][5] , \RF[21][4] , \RF[21][3] , \RF[21][2] ,
         \RF[21][1] , \RF[21][0] , \RF[22][63] , \RF[22][62] , \RF[22][61] ,
         \RF[22][60] , \RF[22][59] , \RF[22][58] , \RF[22][57] , \RF[22][56] ,
         \RF[22][55] , \RF[22][54] , \RF[22][53] , \RF[22][52] , \RF[22][51] ,
         \RF[22][50] , \RF[22][49] , \RF[22][48] , \RF[22][47] , \RF[22][46] ,
         \RF[22][45] , \RF[22][44] , \RF[22][43] , \RF[22][42] , \RF[22][41] ,
         \RF[22][40] , \RF[22][39] , \RF[22][38] , \RF[22][37] , \RF[22][36] ,
         \RF[22][35] , \RF[22][34] , \RF[22][33] , \RF[22][32] , \RF[22][31] ,
         \RF[22][30] , \RF[22][29] , \RF[22][28] , \RF[22][27] , \RF[22][26] ,
         \RF[22][25] , \RF[22][24] , \RF[22][23] , \RF[22][22] , \RF[22][21] ,
         \RF[22][20] , \RF[22][19] , \RF[22][18] , \RF[22][17] , \RF[22][16] ,
         \RF[22][15] , \RF[22][14] , \RF[22][13] , \RF[22][12] , \RF[22][11] ,
         \RF[22][10] , \RF[22][9] , \RF[22][8] , \RF[22][7] , \RF[22][6] ,
         \RF[22][5] , \RF[22][4] , \RF[22][3] , \RF[22][2] , \RF[22][1] ,
         \RF[22][0] , \RF[23][63] , \RF[23][62] , \RF[23][61] , \RF[23][60] ,
         \RF[23][59] , \RF[23][58] , \RF[23][57] , \RF[23][56] , \RF[23][55] ,
         \RF[23][54] , \RF[23][53] , \RF[23][52] , \RF[23][51] , \RF[23][50] ,
         \RF[23][49] , \RF[23][48] , \RF[23][47] , \RF[23][46] , \RF[23][45] ,
         \RF[23][44] , \RF[23][43] , \RF[23][42] , \RF[23][41] , \RF[23][40] ,
         \RF[23][39] , \RF[23][38] , \RF[23][37] , \RF[23][36] , \RF[23][35] ,
         \RF[23][34] , \RF[23][33] , \RF[23][32] , \RF[23][31] , \RF[23][30] ,
         \RF[23][29] , \RF[23][28] , \RF[23][27] , \RF[23][26] , \RF[23][25] ,
         \RF[23][24] , \RF[23][23] , \RF[23][22] , \RF[23][21] , \RF[23][20] ,
         \RF[23][19] , \RF[23][18] , \RF[23][17] , \RF[23][16] , \RF[23][15] ,
         \RF[23][14] , \RF[23][13] , \RF[23][12] , \RF[23][11] , \RF[23][10] ,
         \RF[23][9] , \RF[23][8] , \RF[23][7] , \RF[23][6] , \RF[23][5] ,
         \RF[23][4] , \RF[23][3] , \RF[23][2] , \RF[23][1] , \RF[23][0] ,
         \RF[24][63] , \RF[24][62] , \RF[24][61] , \RF[24][60] , \RF[24][59] ,
         \RF[24][58] , \RF[24][57] , \RF[24][56] , \RF[24][55] , \RF[24][54] ,
         \RF[24][53] , \RF[24][52] , \RF[24][51] , \RF[24][50] , \RF[24][49] ,
         \RF[24][48] , \RF[24][47] , \RF[24][46] , \RF[24][45] , \RF[24][44] ,
         \RF[24][43] , \RF[24][42] , \RF[24][41] , \RF[24][40] , \RF[24][39] ,
         \RF[24][38] , \RF[24][37] , \RF[24][36] , \RF[24][35] , \RF[24][34] ,
         \RF[24][33] , \RF[24][32] , \RF[24][31] , \RF[24][30] , \RF[24][29] ,
         \RF[24][28] , \RF[24][27] , \RF[24][26] , \RF[24][25] , \RF[24][24] ,
         \RF[24][23] , \RF[24][22] , \RF[24][21] , \RF[24][20] , \RF[24][19] ,
         \RF[24][18] , \RF[24][17] , \RF[24][16] , \RF[24][15] , \RF[24][14] ,
         \RF[24][13] , \RF[24][12] , \RF[24][11] , \RF[24][10] , \RF[24][9] ,
         \RF[24][8] , \RF[24][7] , \RF[24][6] , \RF[24][5] , \RF[24][4] ,
         \RF[24][3] , \RF[24][2] , \RF[24][1] , \RF[24][0] , \RF[25][63] ,
         \RF[25][62] , \RF[25][61] , \RF[25][60] , \RF[25][59] , \RF[25][58] ,
         \RF[25][57] , \RF[25][56] , \RF[25][55] , \RF[25][54] , \RF[25][53] ,
         \RF[25][52] , \RF[25][51] , \RF[25][50] , \RF[25][49] , \RF[25][48] ,
         \RF[25][47] , \RF[25][46] , \RF[25][45] , \RF[25][44] , \RF[25][43] ,
         \RF[25][42] , \RF[25][41] , \RF[25][40] , \RF[25][39] , \RF[25][38] ,
         \RF[25][37] , \RF[25][36] , \RF[25][35] , \RF[25][34] , \RF[25][33] ,
         \RF[25][32] , \RF[25][31] , \RF[25][30] , \RF[25][29] , \RF[25][28] ,
         \RF[25][27] , \RF[25][26] , \RF[25][25] , \RF[25][24] , \RF[25][23] ,
         \RF[25][22] , \RF[25][21] , \RF[25][20] , \RF[25][19] , \RF[25][18] ,
         \RF[25][17] , \RF[25][16] , \RF[25][15] , \RF[25][14] , \RF[25][13] ,
         \RF[25][12] , \RF[25][11] , \RF[25][10] , \RF[25][9] , \RF[25][8] ,
         \RF[25][7] , \RF[25][6] , \RF[25][5] , \RF[25][4] , \RF[25][3] ,
         \RF[25][2] , \RF[25][1] , \RF[25][0] , \RF[26][63] , \RF[26][62] ,
         \RF[26][61] , \RF[26][60] , \RF[26][59] , \RF[26][58] , \RF[26][57] ,
         \RF[26][56] , \RF[26][55] , \RF[26][54] , \RF[26][53] , \RF[26][52] ,
         \RF[26][51] , \RF[26][50] , \RF[26][49] , \RF[26][48] , \RF[26][47] ,
         \RF[26][46] , \RF[26][45] , \RF[26][44] , \RF[26][43] , \RF[26][42] ,
         \RF[26][41] , \RF[26][40] , \RF[26][39] , \RF[26][38] , \RF[26][37] ,
         \RF[26][36] , \RF[26][35] , \RF[26][34] , \RF[26][33] , \RF[26][32] ,
         \RF[26][31] , \RF[26][30] , \RF[26][29] , \RF[26][28] , \RF[26][27] ,
         \RF[26][26] , \RF[26][25] , \RF[26][24] , \RF[26][23] , \RF[26][22] ,
         \RF[26][21] , \RF[26][20] , \RF[26][19] , \RF[26][18] , \RF[26][17] ,
         \RF[26][16] , \RF[26][15] , \RF[26][14] , \RF[26][13] , \RF[26][12] ,
         \RF[26][11] , \RF[26][10] , \RF[26][9] , \RF[26][8] , \RF[26][7] ,
         \RF[26][6] , \RF[26][5] , \RF[26][4] , \RF[26][3] , \RF[26][2] ,
         \RF[26][1] , \RF[26][0] , \RF[27][63] , \RF[27][62] , \RF[27][61] ,
         \RF[27][60] , \RF[27][59] , \RF[27][58] , \RF[27][57] , \RF[27][56] ,
         \RF[27][55] , \RF[27][54] , \RF[27][53] , \RF[27][52] , \RF[27][51] ,
         \RF[27][50] , \RF[27][49] , \RF[27][48] , \RF[27][47] , \RF[27][46] ,
         \RF[27][45] , \RF[27][44] , \RF[27][43] , \RF[27][42] , \RF[27][41] ,
         \RF[27][40] , \RF[27][39] , \RF[27][38] , \RF[27][37] , \RF[27][36] ,
         \RF[27][35] , \RF[27][34] , \RF[27][33] , \RF[27][32] , \RF[27][31] ,
         \RF[27][30] , \RF[27][29] , \RF[27][28] , \RF[27][27] , \RF[27][26] ,
         \RF[27][25] , \RF[27][24] , \RF[27][23] , \RF[27][22] , \RF[27][21] ,
         \RF[27][20] , \RF[27][19] , \RF[27][18] , \RF[27][17] , \RF[27][16] ,
         \RF[27][15] , \RF[27][14] , \RF[27][13] , \RF[27][12] , \RF[27][11] ,
         \RF[27][10] , \RF[27][9] , \RF[27][8] , \RF[27][7] , \RF[27][6] ,
         \RF[27][5] , \RF[27][4] , \RF[27][3] , \RF[27][2] , \RF[27][1] ,
         \RF[27][0] , \RF[28][63] , \RF[28][62] , \RF[28][61] , \RF[28][60] ,
         \RF[28][59] , \RF[28][58] , \RF[28][57] , \RF[28][56] , \RF[28][55] ,
         \RF[28][54] , \RF[28][53] , \RF[28][52] , \RF[28][51] , \RF[28][50] ,
         \RF[28][49] , \RF[28][48] , \RF[28][47] , \RF[28][46] , \RF[28][45] ,
         \RF[28][44] , \RF[28][43] , \RF[28][42] , \RF[28][41] , \RF[28][40] ,
         \RF[28][39] , \RF[28][38] , \RF[28][37] , \RF[28][36] , \RF[28][35] ,
         \RF[28][34] , \RF[28][33] , \RF[28][32] , \RF[28][31] , \RF[28][30] ,
         \RF[28][29] , \RF[28][28] , \RF[28][27] , \RF[28][26] , \RF[28][25] ,
         \RF[28][24] , \RF[28][23] , \RF[28][22] , \RF[28][21] , \RF[28][20] ,
         \RF[28][19] , \RF[28][18] , \RF[28][17] , \RF[28][16] , \RF[28][15] ,
         \RF[28][14] , \RF[28][13] , \RF[28][12] , \RF[28][11] , \RF[28][10] ,
         \RF[28][9] , \RF[28][8] , \RF[28][7] , \RF[28][6] , \RF[28][5] ,
         \RF[28][4] , \RF[28][3] , \RF[28][2] , \RF[28][1] , \RF[28][0] ,
         \RF[29][63] , \RF[29][62] , \RF[29][61] , \RF[29][60] , \RF[29][59] ,
         \RF[29][58] , \RF[29][57] , \RF[29][56] , \RF[29][55] , \RF[29][54] ,
         \RF[29][53] , \RF[29][52] , \RF[29][51] , \RF[29][50] , \RF[29][49] ,
         \RF[29][48] , \RF[29][47] , \RF[29][46] , \RF[29][45] , \RF[29][44] ,
         \RF[29][43] , \RF[29][42] , \RF[29][41] , \RF[29][40] , \RF[29][39] ,
         \RF[29][38] , \RF[29][37] , \RF[29][36] , \RF[29][35] , \RF[29][34] ,
         \RF[29][33] , \RF[29][32] , \RF[29][31] , \RF[29][30] , \RF[29][29] ,
         \RF[29][28] , \RF[29][27] , \RF[29][26] , \RF[29][25] , \RF[29][24] ,
         \RF[29][23] , \RF[29][22] , \RF[29][21] , \RF[29][20] , \RF[29][19] ,
         \RF[29][18] , \RF[29][17] , \RF[29][16] , \RF[29][15] , \RF[29][14] ,
         \RF[29][13] , \RF[29][12] , \RF[29][11] , \RF[29][10] , \RF[29][9] ,
         \RF[29][8] , \RF[29][7] , \RF[29][6] , \RF[29][5] , \RF[29][4] ,
         \RF[29][3] , \RF[29][2] , \RF[29][1] , \RF[29][0] , \RF[30][63] ,
         \RF[30][62] , \RF[30][61] , \RF[30][60] , \RF[30][59] , \RF[30][58] ,
         \RF[30][57] , \RF[30][56] , \RF[30][55] , \RF[30][54] , \RF[30][53] ,
         \RF[30][52] , \RF[30][51] , \RF[30][50] , \RF[30][49] , \RF[30][48] ,
         \RF[30][47] , \RF[30][46] , \RF[30][45] , \RF[30][44] , \RF[30][43] ,
         \RF[30][42] , \RF[30][41] , \RF[30][40] , \RF[30][39] , \RF[30][38] ,
         \RF[30][37] , \RF[30][36] , \RF[30][35] , \RF[30][34] , \RF[30][33] ,
         \RF[30][32] , \RF[30][31] , \RF[30][30] , \RF[30][29] , \RF[30][28] ,
         \RF[30][27] , \RF[30][26] , \RF[30][25] , \RF[30][24] , \RF[30][23] ,
         \RF[30][22] , \RF[30][21] , \RF[30][20] , \RF[30][19] , \RF[30][18] ,
         \RF[30][17] , \RF[30][16] , \RF[30][15] , \RF[30][14] , \RF[30][13] ,
         \RF[30][12] , \RF[30][11] , \RF[30][10] , \RF[30][9] , \RF[30][8] ,
         \RF[30][7] , \RF[30][6] , \RF[30][5] , \RF[30][4] , \RF[30][3] ,
         \RF[30][2] , \RF[30][1] , \RF[30][0] , \RF[31][63] , \RF[31][62] ,
         \RF[31][61] , \RF[31][60] , \RF[31][59] , \RF[31][58] , \RF[31][57] ,
         \RF[31][56] , \RF[31][55] , \RF[31][54] , \RF[31][53] , \RF[31][52] ,
         \RF[31][51] , \RF[31][50] , \RF[31][49] , \RF[31][48] , \RF[31][47] ,
         \RF[31][46] , \RF[31][45] , \RF[31][44] , \RF[31][43] , \RF[31][42] ,
         \RF[31][41] , \RF[31][40] , \RF[31][39] , \RF[31][38] , \RF[31][37] ,
         \RF[31][36] , \RF[31][35] , \RF[31][34] , \RF[31][33] , \RF[31][32] ,
         \RF[31][31] , \RF[31][30] , \RF[31][29] , \RF[31][28] , \RF[31][27] ,
         \RF[31][26] , \RF[31][25] , \RF[31][24] , \RF[31][23] , \RF[31][22] ,
         \RF[31][21] , \RF[31][20] , \RF[31][19] , \RF[31][18] , \RF[31][17] ,
         \RF[31][16] , \RF[31][15] , \RF[31][14] , \RF[31][13] , \RF[31][12] ,
         \RF[31][11] , \RF[31][10] , \RF[31][9] , \RF[31][8] , \RF[31][7] ,
         \RF[31][6] , \RF[31][5] , \RF[31][4] , \RF[31][3] , \RF[31][2] ,
         \RF[31][1] , \RF[31][0] , N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74,
         N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N89,
         N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102,
         N103, N104, N105, N106, N107, N108, N109, N110, N111, N112, N113,
         N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, N124,
         N125, N126, N127, N128, N129, N130, N131, N132, N133, N134, N135,
         N136, N137, N138, N139, N140, N141, N142, N143, N144, N145, N146,
         N147, N148, N149, N150, N151, N152, n39, n41, n43, n45, n47, n49, n51,
         n53, n55, n57, n59, n61, n63, n65, n67, n69, n71, n73, n75, n77, n79,
         n81, n83, n85, n87, n89, n91, n93, n95, n97, n99, n101, n103, n105,
         n107, n109, n111, n113, n115, n117, n119, n121, n123, n125, n127,
         n129, n131, n133, n135, n137, n139, n141, n143, n145, n147, n149,
         n151, n153, n155, n157, n159, n161, n163, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835;
  assign N13 = raddr_0[0];
  assign N14 = raddr_0[1];
  assign N15 = raddr_0[2];
  assign N16 = raddr_0[3];
  assign N17 = raddr_0[4];
  assign N18 = raddr_1[0];
  assign N19 = raddr_1[1];
  assign N20 = raddr_1[2];
  assign N21 = raddr_1[3];
  assign N22 = raddr_1[4];

  DFFPOSX1 \RF_reg[0][63]  ( .D(n4242), .CLK(clk), .Q(\RF[0][63] ) );
  DFFPOSX1 \RF_reg[0][62]  ( .D(n4241), .CLK(clk), .Q(\RF[0][62] ) );
  DFFPOSX1 \RF_reg[0][61]  ( .D(n4240), .CLK(clk), .Q(\RF[0][61] ) );
  DFFPOSX1 \RF_reg[0][60]  ( .D(n4239), .CLK(clk), .Q(\RF[0][60] ) );
  DFFPOSX1 \RF_reg[0][59]  ( .D(n4238), .CLK(clk), .Q(\RF[0][59] ) );
  DFFPOSX1 \RF_reg[0][58]  ( .D(n4237), .CLK(clk), .Q(\RF[0][58] ) );
  DFFPOSX1 \RF_reg[0][57]  ( .D(n4236), .CLK(clk), .Q(\RF[0][57] ) );
  DFFPOSX1 \RF_reg[0][56]  ( .D(n4235), .CLK(clk), .Q(\RF[0][56] ) );
  DFFPOSX1 \RF_reg[0][55]  ( .D(n4234), .CLK(clk), .Q(\RF[0][55] ) );
  DFFPOSX1 \RF_reg[0][54]  ( .D(n4233), .CLK(clk), .Q(\RF[0][54] ) );
  DFFPOSX1 \RF_reg[0][53]  ( .D(n4232), .CLK(clk), .Q(\RF[0][53] ) );
  DFFPOSX1 \RF_reg[0][52]  ( .D(n4231), .CLK(clk), .Q(\RF[0][52] ) );
  DFFPOSX1 \RF_reg[0][51]  ( .D(n4230), .CLK(clk), .Q(\RF[0][51] ) );
  DFFPOSX1 \RF_reg[0][50]  ( .D(n4229), .CLK(clk), .Q(\RF[0][50] ) );
  DFFPOSX1 \RF_reg[0][49]  ( .D(n4228), .CLK(clk), .Q(\RF[0][49] ) );
  DFFPOSX1 \RF_reg[0][48]  ( .D(n4227), .CLK(clk), .Q(\RF[0][48] ) );
  DFFPOSX1 \RF_reg[0][47]  ( .D(n4226), .CLK(clk), .Q(\RF[0][47] ) );
  DFFPOSX1 \RF_reg[0][46]  ( .D(n4225), .CLK(clk), .Q(\RF[0][46] ) );
  DFFPOSX1 \RF_reg[0][45]  ( .D(n4224), .CLK(clk), .Q(\RF[0][45] ) );
  DFFPOSX1 \RF_reg[0][44]  ( .D(n4223), .CLK(clk), .Q(\RF[0][44] ) );
  DFFPOSX1 \RF_reg[0][43]  ( .D(n4222), .CLK(clk), .Q(\RF[0][43] ) );
  DFFPOSX1 \RF_reg[0][42]  ( .D(n4221), .CLK(clk), .Q(\RF[0][42] ) );
  DFFPOSX1 \RF_reg[0][41]  ( .D(n4220), .CLK(clk), .Q(\RF[0][41] ) );
  DFFPOSX1 \RF_reg[0][40]  ( .D(n4219), .CLK(clk), .Q(\RF[0][40] ) );
  DFFPOSX1 \RF_reg[0][39]  ( .D(n4218), .CLK(clk), .Q(\RF[0][39] ) );
  DFFPOSX1 \RF_reg[0][38]  ( .D(n4217), .CLK(clk), .Q(\RF[0][38] ) );
  DFFPOSX1 \RF_reg[0][37]  ( .D(n4216), .CLK(clk), .Q(\RF[0][37] ) );
  DFFPOSX1 \RF_reg[0][36]  ( .D(n4215), .CLK(clk), .Q(\RF[0][36] ) );
  DFFPOSX1 \RF_reg[0][35]  ( .D(n4214), .CLK(clk), .Q(\RF[0][35] ) );
  DFFPOSX1 \RF_reg[0][34]  ( .D(n4213), .CLK(clk), .Q(\RF[0][34] ) );
  DFFPOSX1 \RF_reg[0][33]  ( .D(n4212), .CLK(clk), .Q(\RF[0][33] ) );
  DFFPOSX1 \RF_reg[0][32]  ( .D(n4211), .CLK(clk), .Q(\RF[0][32] ) );
  DFFPOSX1 \RF_reg[0][31]  ( .D(n4210), .CLK(clk), .Q(\RF[0][31] ) );
  DFFPOSX1 \RF_reg[0][30]  ( .D(n4209), .CLK(clk), .Q(\RF[0][30] ) );
  DFFPOSX1 \RF_reg[0][29]  ( .D(n4208), .CLK(clk), .Q(\RF[0][29] ) );
  DFFPOSX1 \RF_reg[0][28]  ( .D(n4207), .CLK(clk), .Q(\RF[0][28] ) );
  DFFPOSX1 \RF_reg[0][27]  ( .D(n4206), .CLK(clk), .Q(\RF[0][27] ) );
  DFFPOSX1 \RF_reg[0][26]  ( .D(n4205), .CLK(clk), .Q(\RF[0][26] ) );
  DFFPOSX1 \RF_reg[0][25]  ( .D(n4204), .CLK(clk), .Q(\RF[0][25] ) );
  DFFPOSX1 \RF_reg[0][24]  ( .D(n4203), .CLK(clk), .Q(\RF[0][24] ) );
  DFFPOSX1 \RF_reg[0][23]  ( .D(n4202), .CLK(clk), .Q(\RF[0][23] ) );
  DFFPOSX1 \RF_reg[0][22]  ( .D(n4201), .CLK(clk), .Q(\RF[0][22] ) );
  DFFPOSX1 \RF_reg[0][21]  ( .D(n4200), .CLK(clk), .Q(\RF[0][21] ) );
  DFFPOSX1 \RF_reg[0][20]  ( .D(n4199), .CLK(clk), .Q(\RF[0][20] ) );
  DFFPOSX1 \RF_reg[0][19]  ( .D(n4198), .CLK(clk), .Q(\RF[0][19] ) );
  DFFPOSX1 \RF_reg[0][18]  ( .D(n4197), .CLK(clk), .Q(\RF[0][18] ) );
  DFFPOSX1 \RF_reg[0][17]  ( .D(n4196), .CLK(clk), .Q(\RF[0][17] ) );
  DFFPOSX1 \RF_reg[0][16]  ( .D(n4195), .CLK(clk), .Q(\RF[0][16] ) );
  DFFPOSX1 \RF_reg[0][15]  ( .D(n4194), .CLK(clk), .Q(\RF[0][15] ) );
  DFFPOSX1 \RF_reg[0][14]  ( .D(n4193), .CLK(clk), .Q(\RF[0][14] ) );
  DFFPOSX1 \RF_reg[0][13]  ( .D(n4192), .CLK(clk), .Q(\RF[0][13] ) );
  DFFPOSX1 \RF_reg[0][12]  ( .D(n4191), .CLK(clk), .Q(\RF[0][12] ) );
  DFFPOSX1 \RF_reg[0][11]  ( .D(n4190), .CLK(clk), .Q(\RF[0][11] ) );
  DFFPOSX1 \RF_reg[0][10]  ( .D(n4189), .CLK(clk), .Q(\RF[0][10] ) );
  DFFPOSX1 \RF_reg[0][9]  ( .D(n4188), .CLK(clk), .Q(\RF[0][9] ) );
  DFFPOSX1 \RF_reg[0][8]  ( .D(n4187), .CLK(clk), .Q(\RF[0][8] ) );
  DFFPOSX1 \RF_reg[0][7]  ( .D(n4186), .CLK(clk), .Q(\RF[0][7] ) );
  DFFPOSX1 \RF_reg[0][6]  ( .D(n4185), .CLK(clk), .Q(\RF[0][6] ) );
  DFFPOSX1 \RF_reg[0][5]  ( .D(n4184), .CLK(clk), .Q(\RF[0][5] ) );
  DFFPOSX1 \RF_reg[0][4]  ( .D(n4183), .CLK(clk), .Q(\RF[0][4] ) );
  DFFPOSX1 \RF_reg[0][3]  ( .D(n4182), .CLK(clk), .Q(\RF[0][3] ) );
  DFFPOSX1 \RF_reg[0][2]  ( .D(n4181), .CLK(clk), .Q(\RF[0][2] ) );
  DFFPOSX1 \RF_reg[0][1]  ( .D(n4180), .CLK(clk), .Q(\RF[0][1] ) );
  DFFPOSX1 \RF_reg[0][0]  ( .D(n4179), .CLK(clk), .Q(\RF[0][0] ) );
  DFFPOSX1 \RF_reg[1][63]  ( .D(n4178), .CLK(clk), .Q(\RF[1][63] ) );
  DFFPOSX1 \RF_reg[1][62]  ( .D(n4177), .CLK(clk), .Q(\RF[1][62] ) );
  DFFPOSX1 \RF_reg[1][61]  ( .D(n4176), .CLK(clk), .Q(\RF[1][61] ) );
  DFFPOSX1 \RF_reg[1][60]  ( .D(n4175), .CLK(clk), .Q(\RF[1][60] ) );
  DFFPOSX1 \RF_reg[1][59]  ( .D(n4174), .CLK(clk), .Q(\RF[1][59] ) );
  DFFPOSX1 \RF_reg[1][58]  ( .D(n4173), .CLK(clk), .Q(\RF[1][58] ) );
  DFFPOSX1 \RF_reg[1][57]  ( .D(n4172), .CLK(clk), .Q(\RF[1][57] ) );
  DFFPOSX1 \RF_reg[1][56]  ( .D(n4171), .CLK(clk), .Q(\RF[1][56] ) );
  DFFPOSX1 \RF_reg[1][55]  ( .D(n4170), .CLK(clk), .Q(\RF[1][55] ) );
  DFFPOSX1 \RF_reg[1][54]  ( .D(n4169), .CLK(clk), .Q(\RF[1][54] ) );
  DFFPOSX1 \RF_reg[1][53]  ( .D(n4168), .CLK(clk), .Q(\RF[1][53] ) );
  DFFPOSX1 \RF_reg[1][52]  ( .D(n4167), .CLK(clk), .Q(\RF[1][52] ) );
  DFFPOSX1 \RF_reg[1][51]  ( .D(n4166), .CLK(clk), .Q(\RF[1][51] ) );
  DFFPOSX1 \RF_reg[1][50]  ( .D(n4165), .CLK(clk), .Q(\RF[1][50] ) );
  DFFPOSX1 \RF_reg[1][49]  ( .D(n4164), .CLK(clk), .Q(\RF[1][49] ) );
  DFFPOSX1 \RF_reg[1][48]  ( .D(n4163), .CLK(clk), .Q(\RF[1][48] ) );
  DFFPOSX1 \RF_reg[1][47]  ( .D(n4162), .CLK(clk), .Q(\RF[1][47] ) );
  DFFPOSX1 \RF_reg[1][46]  ( .D(n4161), .CLK(clk), .Q(\RF[1][46] ) );
  DFFPOSX1 \RF_reg[1][45]  ( .D(n4160), .CLK(clk), .Q(\RF[1][45] ) );
  DFFPOSX1 \RF_reg[1][44]  ( .D(n4159), .CLK(clk), .Q(\RF[1][44] ) );
  DFFPOSX1 \RF_reg[1][43]  ( .D(n4158), .CLK(clk), .Q(\RF[1][43] ) );
  DFFPOSX1 \RF_reg[1][42]  ( .D(n4157), .CLK(clk), .Q(\RF[1][42] ) );
  DFFPOSX1 \RF_reg[1][41]  ( .D(n4156), .CLK(clk), .Q(\RF[1][41] ) );
  DFFPOSX1 \RF_reg[1][40]  ( .D(n4155), .CLK(clk), .Q(\RF[1][40] ) );
  DFFPOSX1 \RF_reg[1][39]  ( .D(n4154), .CLK(clk), .Q(\RF[1][39] ) );
  DFFPOSX1 \RF_reg[1][38]  ( .D(n4153), .CLK(clk), .Q(\RF[1][38] ) );
  DFFPOSX1 \RF_reg[1][37]  ( .D(n4152), .CLK(clk), .Q(\RF[1][37] ) );
  DFFPOSX1 \RF_reg[1][36]  ( .D(n4151), .CLK(clk), .Q(\RF[1][36] ) );
  DFFPOSX1 \RF_reg[1][35]  ( .D(n4150), .CLK(clk), .Q(\RF[1][35] ) );
  DFFPOSX1 \RF_reg[1][34]  ( .D(n4149), .CLK(clk), .Q(\RF[1][34] ) );
  DFFPOSX1 \RF_reg[1][33]  ( .D(n4148), .CLK(clk), .Q(\RF[1][33] ) );
  DFFPOSX1 \RF_reg[1][32]  ( .D(n4147), .CLK(clk), .Q(\RF[1][32] ) );
  DFFPOSX1 \RF_reg[1][31]  ( .D(n4146), .CLK(clk), .Q(\RF[1][31] ) );
  DFFPOSX1 \RF_reg[1][30]  ( .D(n4145), .CLK(clk), .Q(\RF[1][30] ) );
  DFFPOSX1 \RF_reg[1][29]  ( .D(n4144), .CLK(clk), .Q(\RF[1][29] ) );
  DFFPOSX1 \RF_reg[1][28]  ( .D(n4143), .CLK(clk), .Q(\RF[1][28] ) );
  DFFPOSX1 \RF_reg[1][27]  ( .D(n4142), .CLK(clk), .Q(\RF[1][27] ) );
  DFFPOSX1 \RF_reg[1][26]  ( .D(n4141), .CLK(clk), .Q(\RF[1][26] ) );
  DFFPOSX1 \RF_reg[1][25]  ( .D(n4140), .CLK(clk), .Q(\RF[1][25] ) );
  DFFPOSX1 \RF_reg[1][24]  ( .D(n4139), .CLK(clk), .Q(\RF[1][24] ) );
  DFFPOSX1 \RF_reg[1][23]  ( .D(n4138), .CLK(clk), .Q(\RF[1][23] ) );
  DFFPOSX1 \RF_reg[1][22]  ( .D(n4137), .CLK(clk), .Q(\RF[1][22] ) );
  DFFPOSX1 \RF_reg[1][21]  ( .D(n4136), .CLK(clk), .Q(\RF[1][21] ) );
  DFFPOSX1 \RF_reg[1][20]  ( .D(n4135), .CLK(clk), .Q(\RF[1][20] ) );
  DFFPOSX1 \RF_reg[1][19]  ( .D(n4134), .CLK(clk), .Q(\RF[1][19] ) );
  DFFPOSX1 \RF_reg[1][18]  ( .D(n4133), .CLK(clk), .Q(\RF[1][18] ) );
  DFFPOSX1 \RF_reg[1][17]  ( .D(n4132), .CLK(clk), .Q(\RF[1][17] ) );
  DFFPOSX1 \RF_reg[1][16]  ( .D(n4131), .CLK(clk), .Q(\RF[1][16] ) );
  DFFPOSX1 \RF_reg[1][15]  ( .D(n4130), .CLK(clk), .Q(\RF[1][15] ) );
  DFFPOSX1 \RF_reg[1][14]  ( .D(n4129), .CLK(clk), .Q(\RF[1][14] ) );
  DFFPOSX1 \RF_reg[1][13]  ( .D(n4128), .CLK(clk), .Q(\RF[1][13] ) );
  DFFPOSX1 \RF_reg[1][12]  ( .D(n4127), .CLK(clk), .Q(\RF[1][12] ) );
  DFFPOSX1 \RF_reg[1][11]  ( .D(n4126), .CLK(clk), .Q(\RF[1][11] ) );
  DFFPOSX1 \RF_reg[1][10]  ( .D(n4125), .CLK(clk), .Q(\RF[1][10] ) );
  DFFPOSX1 \RF_reg[1][9]  ( .D(n4124), .CLK(clk), .Q(\RF[1][9] ) );
  DFFPOSX1 \RF_reg[1][8]  ( .D(n4123), .CLK(clk), .Q(\RF[1][8] ) );
  DFFPOSX1 \RF_reg[1][7]  ( .D(n4122), .CLK(clk), .Q(\RF[1][7] ) );
  DFFPOSX1 \RF_reg[1][6]  ( .D(n4121), .CLK(clk), .Q(\RF[1][6] ) );
  DFFPOSX1 \RF_reg[1][5]  ( .D(n4120), .CLK(clk), .Q(\RF[1][5] ) );
  DFFPOSX1 \RF_reg[1][4]  ( .D(n4119), .CLK(clk), .Q(\RF[1][4] ) );
  DFFPOSX1 \RF_reg[1][3]  ( .D(n4118), .CLK(clk), .Q(\RF[1][3] ) );
  DFFPOSX1 \RF_reg[1][2]  ( .D(n4117), .CLK(clk), .Q(\RF[1][2] ) );
  DFFPOSX1 \RF_reg[1][1]  ( .D(n4116), .CLK(clk), .Q(\RF[1][1] ) );
  DFFPOSX1 \RF_reg[1][0]  ( .D(n4115), .CLK(clk), .Q(\RF[1][0] ) );
  DFFPOSX1 \RF_reg[2][63]  ( .D(n4114), .CLK(clk), .Q(\RF[2][63] ) );
  DFFPOSX1 \RF_reg[2][62]  ( .D(n4113), .CLK(clk), .Q(\RF[2][62] ) );
  DFFPOSX1 \RF_reg[2][61]  ( .D(n4112), .CLK(clk), .Q(\RF[2][61] ) );
  DFFPOSX1 \RF_reg[2][60]  ( .D(n4111), .CLK(clk), .Q(\RF[2][60] ) );
  DFFPOSX1 \RF_reg[2][59]  ( .D(n4110), .CLK(clk), .Q(\RF[2][59] ) );
  DFFPOSX1 \RF_reg[2][58]  ( .D(n4109), .CLK(clk), .Q(\RF[2][58] ) );
  DFFPOSX1 \RF_reg[2][57]  ( .D(n4108), .CLK(clk), .Q(\RF[2][57] ) );
  DFFPOSX1 \RF_reg[2][56]  ( .D(n4107), .CLK(clk), .Q(\RF[2][56] ) );
  DFFPOSX1 \RF_reg[2][55]  ( .D(n4106), .CLK(clk), .Q(\RF[2][55] ) );
  DFFPOSX1 \RF_reg[2][54]  ( .D(n4105), .CLK(clk), .Q(\RF[2][54] ) );
  DFFPOSX1 \RF_reg[2][53]  ( .D(n4104), .CLK(clk), .Q(\RF[2][53] ) );
  DFFPOSX1 \RF_reg[2][52]  ( .D(n4103), .CLK(clk), .Q(\RF[2][52] ) );
  DFFPOSX1 \RF_reg[2][51]  ( .D(n4102), .CLK(clk), .Q(\RF[2][51] ) );
  DFFPOSX1 \RF_reg[2][50]  ( .D(n4101), .CLK(clk), .Q(\RF[2][50] ) );
  DFFPOSX1 \RF_reg[2][49]  ( .D(n4100), .CLK(clk), .Q(\RF[2][49] ) );
  DFFPOSX1 \RF_reg[2][48]  ( .D(n4099), .CLK(clk), .Q(\RF[2][48] ) );
  DFFPOSX1 \RF_reg[2][47]  ( .D(n4098), .CLK(clk), .Q(\RF[2][47] ) );
  DFFPOSX1 \RF_reg[2][46]  ( .D(n4097), .CLK(clk), .Q(\RF[2][46] ) );
  DFFPOSX1 \RF_reg[2][45]  ( .D(n4096), .CLK(clk), .Q(\RF[2][45] ) );
  DFFPOSX1 \RF_reg[2][44]  ( .D(n4095), .CLK(clk), .Q(\RF[2][44] ) );
  DFFPOSX1 \RF_reg[2][43]  ( .D(n4094), .CLK(clk), .Q(\RF[2][43] ) );
  DFFPOSX1 \RF_reg[2][42]  ( .D(n4093), .CLK(clk), .Q(\RF[2][42] ) );
  DFFPOSX1 \RF_reg[2][41]  ( .D(n4092), .CLK(clk), .Q(\RF[2][41] ) );
  DFFPOSX1 \RF_reg[2][40]  ( .D(n4091), .CLK(clk), .Q(\RF[2][40] ) );
  DFFPOSX1 \RF_reg[2][39]  ( .D(n4090), .CLK(clk), .Q(\RF[2][39] ) );
  DFFPOSX1 \RF_reg[2][38]  ( .D(n4089), .CLK(clk), .Q(\RF[2][38] ) );
  DFFPOSX1 \RF_reg[2][37]  ( .D(n4088), .CLK(clk), .Q(\RF[2][37] ) );
  DFFPOSX1 \RF_reg[2][36]  ( .D(n4087), .CLK(clk), .Q(\RF[2][36] ) );
  DFFPOSX1 \RF_reg[2][35]  ( .D(n4086), .CLK(clk), .Q(\RF[2][35] ) );
  DFFPOSX1 \RF_reg[2][34]  ( .D(n4085), .CLK(clk), .Q(\RF[2][34] ) );
  DFFPOSX1 \RF_reg[2][33]  ( .D(n4084), .CLK(clk), .Q(\RF[2][33] ) );
  DFFPOSX1 \RF_reg[2][32]  ( .D(n4083), .CLK(clk), .Q(\RF[2][32] ) );
  DFFPOSX1 \RF_reg[2][31]  ( .D(n4082), .CLK(clk), .Q(\RF[2][31] ) );
  DFFPOSX1 \RF_reg[2][30]  ( .D(n4081), .CLK(clk), .Q(\RF[2][30] ) );
  DFFPOSX1 \RF_reg[2][29]  ( .D(n4080), .CLK(clk), .Q(\RF[2][29] ) );
  DFFPOSX1 \RF_reg[2][28]  ( .D(n4079), .CLK(clk), .Q(\RF[2][28] ) );
  DFFPOSX1 \RF_reg[2][27]  ( .D(n4078), .CLK(clk), .Q(\RF[2][27] ) );
  DFFPOSX1 \RF_reg[2][26]  ( .D(n4077), .CLK(clk), .Q(\RF[2][26] ) );
  DFFPOSX1 \RF_reg[2][25]  ( .D(n4076), .CLK(clk), .Q(\RF[2][25] ) );
  DFFPOSX1 \RF_reg[2][24]  ( .D(n4075), .CLK(clk), .Q(\RF[2][24] ) );
  DFFPOSX1 \RF_reg[2][23]  ( .D(n4074), .CLK(clk), .Q(\RF[2][23] ) );
  DFFPOSX1 \RF_reg[2][22]  ( .D(n4073), .CLK(clk), .Q(\RF[2][22] ) );
  DFFPOSX1 \RF_reg[2][21]  ( .D(n4072), .CLK(clk), .Q(\RF[2][21] ) );
  DFFPOSX1 \RF_reg[2][20]  ( .D(n4071), .CLK(clk), .Q(\RF[2][20] ) );
  DFFPOSX1 \RF_reg[2][19]  ( .D(n4070), .CLK(clk), .Q(\RF[2][19] ) );
  DFFPOSX1 \RF_reg[2][18]  ( .D(n4069), .CLK(clk), .Q(\RF[2][18] ) );
  DFFPOSX1 \RF_reg[2][17]  ( .D(n4068), .CLK(clk), .Q(\RF[2][17] ) );
  DFFPOSX1 \RF_reg[2][16]  ( .D(n4067), .CLK(clk), .Q(\RF[2][16] ) );
  DFFPOSX1 \RF_reg[2][15]  ( .D(n4066), .CLK(clk), .Q(\RF[2][15] ) );
  DFFPOSX1 \RF_reg[2][14]  ( .D(n4065), .CLK(clk), .Q(\RF[2][14] ) );
  DFFPOSX1 \RF_reg[2][13]  ( .D(n4064), .CLK(clk), .Q(\RF[2][13] ) );
  DFFPOSX1 \RF_reg[2][12]  ( .D(n4063), .CLK(clk), .Q(\RF[2][12] ) );
  DFFPOSX1 \RF_reg[2][11]  ( .D(n4062), .CLK(clk), .Q(\RF[2][11] ) );
  DFFPOSX1 \RF_reg[2][10]  ( .D(n4061), .CLK(clk), .Q(\RF[2][10] ) );
  DFFPOSX1 \RF_reg[2][9]  ( .D(n4060), .CLK(clk), .Q(\RF[2][9] ) );
  DFFPOSX1 \RF_reg[2][8]  ( .D(n4059), .CLK(clk), .Q(\RF[2][8] ) );
  DFFPOSX1 \RF_reg[2][7]  ( .D(n4058), .CLK(clk), .Q(\RF[2][7] ) );
  DFFPOSX1 \RF_reg[2][6]  ( .D(n4057), .CLK(clk), .Q(\RF[2][6] ) );
  DFFPOSX1 \RF_reg[2][5]  ( .D(n4056), .CLK(clk), .Q(\RF[2][5] ) );
  DFFPOSX1 \RF_reg[2][4]  ( .D(n4055), .CLK(clk), .Q(\RF[2][4] ) );
  DFFPOSX1 \RF_reg[2][3]  ( .D(n4054), .CLK(clk), .Q(\RF[2][3] ) );
  DFFPOSX1 \RF_reg[2][2]  ( .D(n4053), .CLK(clk), .Q(\RF[2][2] ) );
  DFFPOSX1 \RF_reg[2][1]  ( .D(n4052), .CLK(clk), .Q(\RF[2][1] ) );
  DFFPOSX1 \RF_reg[2][0]  ( .D(n4051), .CLK(clk), .Q(\RF[2][0] ) );
  DFFPOSX1 \RF_reg[3][63]  ( .D(n4050), .CLK(clk), .Q(\RF[3][63] ) );
  DFFPOSX1 \RF_reg[3][62]  ( .D(n4049), .CLK(clk), .Q(\RF[3][62] ) );
  DFFPOSX1 \RF_reg[3][61]  ( .D(n4048), .CLK(clk), .Q(\RF[3][61] ) );
  DFFPOSX1 \RF_reg[3][60]  ( .D(n4047), .CLK(clk), .Q(\RF[3][60] ) );
  DFFPOSX1 \RF_reg[3][59]  ( .D(n4046), .CLK(clk), .Q(\RF[3][59] ) );
  DFFPOSX1 \RF_reg[3][58]  ( .D(n4045), .CLK(clk), .Q(\RF[3][58] ) );
  DFFPOSX1 \RF_reg[3][57]  ( .D(n4044), .CLK(clk), .Q(\RF[3][57] ) );
  DFFPOSX1 \RF_reg[3][56]  ( .D(n4043), .CLK(clk), .Q(\RF[3][56] ) );
  DFFPOSX1 \RF_reg[3][55]  ( .D(n4042), .CLK(clk), .Q(\RF[3][55] ) );
  DFFPOSX1 \RF_reg[3][54]  ( .D(n4041), .CLK(clk), .Q(\RF[3][54] ) );
  DFFPOSX1 \RF_reg[3][53]  ( .D(n4040), .CLK(clk), .Q(\RF[3][53] ) );
  DFFPOSX1 \RF_reg[3][52]  ( .D(n4039), .CLK(clk), .Q(\RF[3][52] ) );
  DFFPOSX1 \RF_reg[3][51]  ( .D(n4038), .CLK(clk), .Q(\RF[3][51] ) );
  DFFPOSX1 \RF_reg[3][50]  ( .D(n4037), .CLK(clk), .Q(\RF[3][50] ) );
  DFFPOSX1 \RF_reg[3][49]  ( .D(n4036), .CLK(clk), .Q(\RF[3][49] ) );
  DFFPOSX1 \RF_reg[3][48]  ( .D(n4035), .CLK(clk), .Q(\RF[3][48] ) );
  DFFPOSX1 \RF_reg[3][47]  ( .D(n4034), .CLK(clk), .Q(\RF[3][47] ) );
  DFFPOSX1 \RF_reg[3][46]  ( .D(n4033), .CLK(clk), .Q(\RF[3][46] ) );
  DFFPOSX1 \RF_reg[3][45]  ( .D(n4032), .CLK(clk), .Q(\RF[3][45] ) );
  DFFPOSX1 \RF_reg[3][44]  ( .D(n4031), .CLK(clk), .Q(\RF[3][44] ) );
  DFFPOSX1 \RF_reg[3][43]  ( .D(n4030), .CLK(clk), .Q(\RF[3][43] ) );
  DFFPOSX1 \RF_reg[3][42]  ( .D(n4029), .CLK(clk), .Q(\RF[3][42] ) );
  DFFPOSX1 \RF_reg[3][41]  ( .D(n4028), .CLK(clk), .Q(\RF[3][41] ) );
  DFFPOSX1 \RF_reg[3][40]  ( .D(n4027), .CLK(clk), .Q(\RF[3][40] ) );
  DFFPOSX1 \RF_reg[3][39]  ( .D(n4026), .CLK(clk), .Q(\RF[3][39] ) );
  DFFPOSX1 \RF_reg[3][38]  ( .D(n4025), .CLK(clk), .Q(\RF[3][38] ) );
  DFFPOSX1 \RF_reg[3][37]  ( .D(n4024), .CLK(clk), .Q(\RF[3][37] ) );
  DFFPOSX1 \RF_reg[3][36]  ( .D(n4023), .CLK(clk), .Q(\RF[3][36] ) );
  DFFPOSX1 \RF_reg[3][35]  ( .D(n4022), .CLK(clk), .Q(\RF[3][35] ) );
  DFFPOSX1 \RF_reg[3][34]  ( .D(n4021), .CLK(clk), .Q(\RF[3][34] ) );
  DFFPOSX1 \RF_reg[3][33]  ( .D(n4020), .CLK(clk), .Q(\RF[3][33] ) );
  DFFPOSX1 \RF_reg[3][32]  ( .D(n4019), .CLK(clk), .Q(\RF[3][32] ) );
  DFFPOSX1 \RF_reg[3][31]  ( .D(n4018), .CLK(clk), .Q(\RF[3][31] ) );
  DFFPOSX1 \RF_reg[3][30]  ( .D(n4017), .CLK(clk), .Q(\RF[3][30] ) );
  DFFPOSX1 \RF_reg[3][29]  ( .D(n4016), .CLK(clk), .Q(\RF[3][29] ) );
  DFFPOSX1 \RF_reg[3][28]  ( .D(n4015), .CLK(clk), .Q(\RF[3][28] ) );
  DFFPOSX1 \RF_reg[3][27]  ( .D(n4014), .CLK(clk), .Q(\RF[3][27] ) );
  DFFPOSX1 \RF_reg[3][26]  ( .D(n4013), .CLK(clk), .Q(\RF[3][26] ) );
  DFFPOSX1 \RF_reg[3][25]  ( .D(n4012), .CLK(clk), .Q(\RF[3][25] ) );
  DFFPOSX1 \RF_reg[3][24]  ( .D(n4011), .CLK(clk), .Q(\RF[3][24] ) );
  DFFPOSX1 \RF_reg[3][23]  ( .D(n4010), .CLK(clk), .Q(\RF[3][23] ) );
  DFFPOSX1 \RF_reg[3][22]  ( .D(n4009), .CLK(clk), .Q(\RF[3][22] ) );
  DFFPOSX1 \RF_reg[3][21]  ( .D(n4008), .CLK(clk), .Q(\RF[3][21] ) );
  DFFPOSX1 \RF_reg[3][20]  ( .D(n4007), .CLK(clk), .Q(\RF[3][20] ) );
  DFFPOSX1 \RF_reg[3][19]  ( .D(n4006), .CLK(clk), .Q(\RF[3][19] ) );
  DFFPOSX1 \RF_reg[3][18]  ( .D(n4005), .CLK(clk), .Q(\RF[3][18] ) );
  DFFPOSX1 \RF_reg[3][17]  ( .D(n4004), .CLK(clk), .Q(\RF[3][17] ) );
  DFFPOSX1 \RF_reg[3][16]  ( .D(n4003), .CLK(clk), .Q(\RF[3][16] ) );
  DFFPOSX1 \RF_reg[3][15]  ( .D(n4002), .CLK(clk), .Q(\RF[3][15] ) );
  DFFPOSX1 \RF_reg[3][14]  ( .D(n4001), .CLK(clk), .Q(\RF[3][14] ) );
  DFFPOSX1 \RF_reg[3][13]  ( .D(n4000), .CLK(clk), .Q(\RF[3][13] ) );
  DFFPOSX1 \RF_reg[3][12]  ( .D(n3999), .CLK(clk), .Q(\RF[3][12] ) );
  DFFPOSX1 \RF_reg[3][11]  ( .D(n3998), .CLK(clk), .Q(\RF[3][11] ) );
  DFFPOSX1 \RF_reg[3][10]  ( .D(n3997), .CLK(clk), .Q(\RF[3][10] ) );
  DFFPOSX1 \RF_reg[3][9]  ( .D(n3996), .CLK(clk), .Q(\RF[3][9] ) );
  DFFPOSX1 \RF_reg[3][8]  ( .D(n3995), .CLK(clk), .Q(\RF[3][8] ) );
  DFFPOSX1 \RF_reg[3][7]  ( .D(n3994), .CLK(clk), .Q(\RF[3][7] ) );
  DFFPOSX1 \RF_reg[3][6]  ( .D(n3993), .CLK(clk), .Q(\RF[3][6] ) );
  DFFPOSX1 \RF_reg[3][5]  ( .D(n3992), .CLK(clk), .Q(\RF[3][5] ) );
  DFFPOSX1 \RF_reg[3][4]  ( .D(n3991), .CLK(clk), .Q(\RF[3][4] ) );
  DFFPOSX1 \RF_reg[3][3]  ( .D(n3990), .CLK(clk), .Q(\RF[3][3] ) );
  DFFPOSX1 \RF_reg[3][2]  ( .D(n3989), .CLK(clk), .Q(\RF[3][2] ) );
  DFFPOSX1 \RF_reg[3][1]  ( .D(n3988), .CLK(clk), .Q(\RF[3][1] ) );
  DFFPOSX1 \RF_reg[3][0]  ( .D(n3987), .CLK(clk), .Q(\RF[3][0] ) );
  DFFPOSX1 \RF_reg[4][63]  ( .D(n3986), .CLK(clk), .Q(\RF[4][63] ) );
  DFFPOSX1 \RF_reg[4][62]  ( .D(n3985), .CLK(clk), .Q(\RF[4][62] ) );
  DFFPOSX1 \RF_reg[4][61]  ( .D(n3984), .CLK(clk), .Q(\RF[4][61] ) );
  DFFPOSX1 \RF_reg[4][60]  ( .D(n3983), .CLK(clk), .Q(\RF[4][60] ) );
  DFFPOSX1 \RF_reg[4][59]  ( .D(n3982), .CLK(clk), .Q(\RF[4][59] ) );
  DFFPOSX1 \RF_reg[4][58]  ( .D(n3981), .CLK(clk), .Q(\RF[4][58] ) );
  DFFPOSX1 \RF_reg[4][57]  ( .D(n3980), .CLK(clk), .Q(\RF[4][57] ) );
  DFFPOSX1 \RF_reg[4][56]  ( .D(n3979), .CLK(clk), .Q(\RF[4][56] ) );
  DFFPOSX1 \RF_reg[4][55]  ( .D(n3978), .CLK(clk), .Q(\RF[4][55] ) );
  DFFPOSX1 \RF_reg[4][54]  ( .D(n3977), .CLK(clk), .Q(\RF[4][54] ) );
  DFFPOSX1 \RF_reg[4][53]  ( .D(n3976), .CLK(clk), .Q(\RF[4][53] ) );
  DFFPOSX1 \RF_reg[4][52]  ( .D(n3975), .CLK(clk), .Q(\RF[4][52] ) );
  DFFPOSX1 \RF_reg[4][51]  ( .D(n3974), .CLK(clk), .Q(\RF[4][51] ) );
  DFFPOSX1 \RF_reg[4][50]  ( .D(n3973), .CLK(clk), .Q(\RF[4][50] ) );
  DFFPOSX1 \RF_reg[4][49]  ( .D(n3972), .CLK(clk), .Q(\RF[4][49] ) );
  DFFPOSX1 \RF_reg[4][48]  ( .D(n3971), .CLK(clk), .Q(\RF[4][48] ) );
  DFFPOSX1 \RF_reg[4][47]  ( .D(n3970), .CLK(clk), .Q(\RF[4][47] ) );
  DFFPOSX1 \RF_reg[4][46]  ( .D(n3969), .CLK(clk), .Q(\RF[4][46] ) );
  DFFPOSX1 \RF_reg[4][45]  ( .D(n3968), .CLK(clk), .Q(\RF[4][45] ) );
  DFFPOSX1 \RF_reg[4][44]  ( .D(n3967), .CLK(clk), .Q(\RF[4][44] ) );
  DFFPOSX1 \RF_reg[4][43]  ( .D(n3966), .CLK(clk), .Q(\RF[4][43] ) );
  DFFPOSX1 \RF_reg[4][42]  ( .D(n3965), .CLK(clk), .Q(\RF[4][42] ) );
  DFFPOSX1 \RF_reg[4][41]  ( .D(n3964), .CLK(clk), .Q(\RF[4][41] ) );
  DFFPOSX1 \RF_reg[4][40]  ( .D(n3963), .CLK(clk), .Q(\RF[4][40] ) );
  DFFPOSX1 \RF_reg[4][39]  ( .D(n3962), .CLK(clk), .Q(\RF[4][39] ) );
  DFFPOSX1 \RF_reg[4][38]  ( .D(n3961), .CLK(clk), .Q(\RF[4][38] ) );
  DFFPOSX1 \RF_reg[4][37]  ( .D(n3960), .CLK(clk), .Q(\RF[4][37] ) );
  DFFPOSX1 \RF_reg[4][36]  ( .D(n3959), .CLK(clk), .Q(\RF[4][36] ) );
  DFFPOSX1 \RF_reg[4][35]  ( .D(n3958), .CLK(clk), .Q(\RF[4][35] ) );
  DFFPOSX1 \RF_reg[4][34]  ( .D(n3957), .CLK(clk), .Q(\RF[4][34] ) );
  DFFPOSX1 \RF_reg[4][33]  ( .D(n3956), .CLK(clk), .Q(\RF[4][33] ) );
  DFFPOSX1 \RF_reg[4][32]  ( .D(n3955), .CLK(clk), .Q(\RF[4][32] ) );
  DFFPOSX1 \RF_reg[4][31]  ( .D(n3954), .CLK(clk), .Q(\RF[4][31] ) );
  DFFPOSX1 \RF_reg[4][30]  ( .D(n3953), .CLK(clk), .Q(\RF[4][30] ) );
  DFFPOSX1 \RF_reg[4][29]  ( .D(n3952), .CLK(clk), .Q(\RF[4][29] ) );
  DFFPOSX1 \RF_reg[4][28]  ( .D(n3951), .CLK(clk), .Q(\RF[4][28] ) );
  DFFPOSX1 \RF_reg[4][27]  ( .D(n3950), .CLK(clk), .Q(\RF[4][27] ) );
  DFFPOSX1 \RF_reg[4][26]  ( .D(n3949), .CLK(clk), .Q(\RF[4][26] ) );
  DFFPOSX1 \RF_reg[4][25]  ( .D(n3948), .CLK(clk), .Q(\RF[4][25] ) );
  DFFPOSX1 \RF_reg[4][24]  ( .D(n3947), .CLK(clk), .Q(\RF[4][24] ) );
  DFFPOSX1 \RF_reg[4][23]  ( .D(n3946), .CLK(clk), .Q(\RF[4][23] ) );
  DFFPOSX1 \RF_reg[4][22]  ( .D(n3945), .CLK(clk), .Q(\RF[4][22] ) );
  DFFPOSX1 \RF_reg[4][21]  ( .D(n3944), .CLK(clk), .Q(\RF[4][21] ) );
  DFFPOSX1 \RF_reg[4][20]  ( .D(n3943), .CLK(clk), .Q(\RF[4][20] ) );
  DFFPOSX1 \RF_reg[4][19]  ( .D(n3942), .CLK(clk), .Q(\RF[4][19] ) );
  DFFPOSX1 \RF_reg[4][18]  ( .D(n3941), .CLK(clk), .Q(\RF[4][18] ) );
  DFFPOSX1 \RF_reg[4][17]  ( .D(n3940), .CLK(clk), .Q(\RF[4][17] ) );
  DFFPOSX1 \RF_reg[4][16]  ( .D(n3939), .CLK(clk), .Q(\RF[4][16] ) );
  DFFPOSX1 \RF_reg[4][15]  ( .D(n3938), .CLK(clk), .Q(\RF[4][15] ) );
  DFFPOSX1 \RF_reg[4][14]  ( .D(n3937), .CLK(clk), .Q(\RF[4][14] ) );
  DFFPOSX1 \RF_reg[4][13]  ( .D(n3936), .CLK(clk), .Q(\RF[4][13] ) );
  DFFPOSX1 \RF_reg[4][12]  ( .D(n3935), .CLK(clk), .Q(\RF[4][12] ) );
  DFFPOSX1 \RF_reg[4][11]  ( .D(n3934), .CLK(clk), .Q(\RF[4][11] ) );
  DFFPOSX1 \RF_reg[4][10]  ( .D(n3933), .CLK(clk), .Q(\RF[4][10] ) );
  DFFPOSX1 \RF_reg[4][9]  ( .D(n3932), .CLK(clk), .Q(\RF[4][9] ) );
  DFFPOSX1 \RF_reg[4][8]  ( .D(n3931), .CLK(clk), .Q(\RF[4][8] ) );
  DFFPOSX1 \RF_reg[4][7]  ( .D(n3930), .CLK(clk), .Q(\RF[4][7] ) );
  DFFPOSX1 \RF_reg[4][6]  ( .D(n3929), .CLK(clk), .Q(\RF[4][6] ) );
  DFFPOSX1 \RF_reg[4][5]  ( .D(n3928), .CLK(clk), .Q(\RF[4][5] ) );
  DFFPOSX1 \RF_reg[4][4]  ( .D(n3927), .CLK(clk), .Q(\RF[4][4] ) );
  DFFPOSX1 \RF_reg[4][3]  ( .D(n3926), .CLK(clk), .Q(\RF[4][3] ) );
  DFFPOSX1 \RF_reg[4][2]  ( .D(n3925), .CLK(clk), .Q(\RF[4][2] ) );
  DFFPOSX1 \RF_reg[4][1]  ( .D(n3924), .CLK(clk), .Q(\RF[4][1] ) );
  DFFPOSX1 \RF_reg[4][0]  ( .D(n3923), .CLK(clk), .Q(\RF[4][0] ) );
  DFFPOSX1 \RF_reg[5][63]  ( .D(n3922), .CLK(clk), .Q(\RF[5][63] ) );
  DFFPOSX1 \RF_reg[5][62]  ( .D(n3921), .CLK(clk), .Q(\RF[5][62] ) );
  DFFPOSX1 \RF_reg[5][61]  ( .D(n3920), .CLK(clk), .Q(\RF[5][61] ) );
  DFFPOSX1 \RF_reg[5][60]  ( .D(n3919), .CLK(clk), .Q(\RF[5][60] ) );
  DFFPOSX1 \RF_reg[5][59]  ( .D(n3918), .CLK(clk), .Q(\RF[5][59] ) );
  DFFPOSX1 \RF_reg[5][58]  ( .D(n3917), .CLK(clk), .Q(\RF[5][58] ) );
  DFFPOSX1 \RF_reg[5][57]  ( .D(n3916), .CLK(clk), .Q(\RF[5][57] ) );
  DFFPOSX1 \RF_reg[5][56]  ( .D(n3915), .CLK(clk), .Q(\RF[5][56] ) );
  DFFPOSX1 \RF_reg[5][55]  ( .D(n3914), .CLK(clk), .Q(\RF[5][55] ) );
  DFFPOSX1 \RF_reg[5][54]  ( .D(n3913), .CLK(clk), .Q(\RF[5][54] ) );
  DFFPOSX1 \RF_reg[5][53]  ( .D(n3912), .CLK(clk), .Q(\RF[5][53] ) );
  DFFPOSX1 \RF_reg[5][52]  ( .D(n3911), .CLK(clk), .Q(\RF[5][52] ) );
  DFFPOSX1 \RF_reg[5][51]  ( .D(n3910), .CLK(clk), .Q(\RF[5][51] ) );
  DFFPOSX1 \RF_reg[5][50]  ( .D(n3909), .CLK(clk), .Q(\RF[5][50] ) );
  DFFPOSX1 \RF_reg[5][49]  ( .D(n3908), .CLK(clk), .Q(\RF[5][49] ) );
  DFFPOSX1 \RF_reg[5][48]  ( .D(n3907), .CLK(clk), .Q(\RF[5][48] ) );
  DFFPOSX1 \RF_reg[5][47]  ( .D(n3906), .CLK(clk), .Q(\RF[5][47] ) );
  DFFPOSX1 \RF_reg[5][46]  ( .D(n3905), .CLK(clk), .Q(\RF[5][46] ) );
  DFFPOSX1 \RF_reg[5][45]  ( .D(n3904), .CLK(clk), .Q(\RF[5][45] ) );
  DFFPOSX1 \RF_reg[5][44]  ( .D(n3903), .CLK(clk), .Q(\RF[5][44] ) );
  DFFPOSX1 \RF_reg[5][43]  ( .D(n3902), .CLK(clk), .Q(\RF[5][43] ) );
  DFFPOSX1 \RF_reg[5][42]  ( .D(n3901), .CLK(clk), .Q(\RF[5][42] ) );
  DFFPOSX1 \RF_reg[5][41]  ( .D(n3900), .CLK(clk), .Q(\RF[5][41] ) );
  DFFPOSX1 \RF_reg[5][40]  ( .D(n3899), .CLK(clk), .Q(\RF[5][40] ) );
  DFFPOSX1 \RF_reg[5][39]  ( .D(n3898), .CLK(clk), .Q(\RF[5][39] ) );
  DFFPOSX1 \RF_reg[5][38]  ( .D(n3897), .CLK(clk), .Q(\RF[5][38] ) );
  DFFPOSX1 \RF_reg[5][37]  ( .D(n3896), .CLK(clk), .Q(\RF[5][37] ) );
  DFFPOSX1 \RF_reg[5][36]  ( .D(n3895), .CLK(clk), .Q(\RF[5][36] ) );
  DFFPOSX1 \RF_reg[5][35]  ( .D(n3894), .CLK(clk), .Q(\RF[5][35] ) );
  DFFPOSX1 \RF_reg[5][34]  ( .D(n3893), .CLK(clk), .Q(\RF[5][34] ) );
  DFFPOSX1 \RF_reg[5][33]  ( .D(n3892), .CLK(clk), .Q(\RF[5][33] ) );
  DFFPOSX1 \RF_reg[5][32]  ( .D(n3891), .CLK(clk), .Q(\RF[5][32] ) );
  DFFPOSX1 \RF_reg[5][31]  ( .D(n3890), .CLK(clk), .Q(\RF[5][31] ) );
  DFFPOSX1 \RF_reg[5][30]  ( .D(n3889), .CLK(clk), .Q(\RF[5][30] ) );
  DFFPOSX1 \RF_reg[5][29]  ( .D(n3888), .CLK(clk), .Q(\RF[5][29] ) );
  DFFPOSX1 \RF_reg[5][28]  ( .D(n3887), .CLK(clk), .Q(\RF[5][28] ) );
  DFFPOSX1 \RF_reg[5][27]  ( .D(n3886), .CLK(clk), .Q(\RF[5][27] ) );
  DFFPOSX1 \RF_reg[5][26]  ( .D(n3885), .CLK(clk), .Q(\RF[5][26] ) );
  DFFPOSX1 \RF_reg[5][25]  ( .D(n3884), .CLK(clk), .Q(\RF[5][25] ) );
  DFFPOSX1 \RF_reg[5][24]  ( .D(n3883), .CLK(clk), .Q(\RF[5][24] ) );
  DFFPOSX1 \RF_reg[5][23]  ( .D(n3882), .CLK(clk), .Q(\RF[5][23] ) );
  DFFPOSX1 \RF_reg[5][22]  ( .D(n3881), .CLK(clk), .Q(\RF[5][22] ) );
  DFFPOSX1 \RF_reg[5][21]  ( .D(n3880), .CLK(clk), .Q(\RF[5][21] ) );
  DFFPOSX1 \RF_reg[5][20]  ( .D(n3879), .CLK(clk), .Q(\RF[5][20] ) );
  DFFPOSX1 \RF_reg[5][19]  ( .D(n3878), .CLK(clk), .Q(\RF[5][19] ) );
  DFFPOSX1 \RF_reg[5][18]  ( .D(n3877), .CLK(clk), .Q(\RF[5][18] ) );
  DFFPOSX1 \RF_reg[5][17]  ( .D(n3876), .CLK(clk), .Q(\RF[5][17] ) );
  DFFPOSX1 \RF_reg[5][16]  ( .D(n3875), .CLK(clk), .Q(\RF[5][16] ) );
  DFFPOSX1 \RF_reg[5][15]  ( .D(n3874), .CLK(clk), .Q(\RF[5][15] ) );
  DFFPOSX1 \RF_reg[5][14]  ( .D(n3873), .CLK(clk), .Q(\RF[5][14] ) );
  DFFPOSX1 \RF_reg[5][13]  ( .D(n3872), .CLK(clk), .Q(\RF[5][13] ) );
  DFFPOSX1 \RF_reg[5][12]  ( .D(n3871), .CLK(clk), .Q(\RF[5][12] ) );
  DFFPOSX1 \RF_reg[5][11]  ( .D(n3870), .CLK(clk), .Q(\RF[5][11] ) );
  DFFPOSX1 \RF_reg[5][10]  ( .D(n3869), .CLK(clk), .Q(\RF[5][10] ) );
  DFFPOSX1 \RF_reg[5][9]  ( .D(n3868), .CLK(clk), .Q(\RF[5][9] ) );
  DFFPOSX1 \RF_reg[5][8]  ( .D(n3867), .CLK(clk), .Q(\RF[5][8] ) );
  DFFPOSX1 \RF_reg[5][7]  ( .D(n3866), .CLK(clk), .Q(\RF[5][7] ) );
  DFFPOSX1 \RF_reg[5][6]  ( .D(n3865), .CLK(clk), .Q(\RF[5][6] ) );
  DFFPOSX1 \RF_reg[5][5]  ( .D(n3864), .CLK(clk), .Q(\RF[5][5] ) );
  DFFPOSX1 \RF_reg[5][4]  ( .D(n3863), .CLK(clk), .Q(\RF[5][4] ) );
  DFFPOSX1 \RF_reg[5][3]  ( .D(n3862), .CLK(clk), .Q(\RF[5][3] ) );
  DFFPOSX1 \RF_reg[5][2]  ( .D(n3861), .CLK(clk), .Q(\RF[5][2] ) );
  DFFPOSX1 \RF_reg[5][1]  ( .D(n3860), .CLK(clk), .Q(\RF[5][1] ) );
  DFFPOSX1 \RF_reg[5][0]  ( .D(n3859), .CLK(clk), .Q(\RF[5][0] ) );
  DFFPOSX1 \RF_reg[6][63]  ( .D(n3858), .CLK(clk), .Q(\RF[6][63] ) );
  DFFPOSX1 \RF_reg[6][62]  ( .D(n3857), .CLK(clk), .Q(\RF[6][62] ) );
  DFFPOSX1 \RF_reg[6][61]  ( .D(n3856), .CLK(clk), .Q(\RF[6][61] ) );
  DFFPOSX1 \RF_reg[6][60]  ( .D(n3855), .CLK(clk), .Q(\RF[6][60] ) );
  DFFPOSX1 \RF_reg[6][59]  ( .D(n3854), .CLK(clk), .Q(\RF[6][59] ) );
  DFFPOSX1 \RF_reg[6][58]  ( .D(n3853), .CLK(clk), .Q(\RF[6][58] ) );
  DFFPOSX1 \RF_reg[6][57]  ( .D(n3852), .CLK(clk), .Q(\RF[6][57] ) );
  DFFPOSX1 \RF_reg[6][56]  ( .D(n3851), .CLK(clk), .Q(\RF[6][56] ) );
  DFFPOSX1 \RF_reg[6][55]  ( .D(n3850), .CLK(clk), .Q(\RF[6][55] ) );
  DFFPOSX1 \RF_reg[6][54]  ( .D(n3849), .CLK(clk), .Q(\RF[6][54] ) );
  DFFPOSX1 \RF_reg[6][53]  ( .D(n3848), .CLK(clk), .Q(\RF[6][53] ) );
  DFFPOSX1 \RF_reg[6][52]  ( .D(n3847), .CLK(clk), .Q(\RF[6][52] ) );
  DFFPOSX1 \RF_reg[6][51]  ( .D(n3846), .CLK(clk), .Q(\RF[6][51] ) );
  DFFPOSX1 \RF_reg[6][50]  ( .D(n3845), .CLK(clk), .Q(\RF[6][50] ) );
  DFFPOSX1 \RF_reg[6][49]  ( .D(n3844), .CLK(clk), .Q(\RF[6][49] ) );
  DFFPOSX1 \RF_reg[6][48]  ( .D(n3843), .CLK(clk), .Q(\RF[6][48] ) );
  DFFPOSX1 \RF_reg[6][47]  ( .D(n3842), .CLK(clk), .Q(\RF[6][47] ) );
  DFFPOSX1 \RF_reg[6][46]  ( .D(n3841), .CLK(clk), .Q(\RF[6][46] ) );
  DFFPOSX1 \RF_reg[6][45]  ( .D(n3840), .CLK(clk), .Q(\RF[6][45] ) );
  DFFPOSX1 \RF_reg[6][44]  ( .D(n3839), .CLK(clk), .Q(\RF[6][44] ) );
  DFFPOSX1 \RF_reg[6][43]  ( .D(n3838), .CLK(clk), .Q(\RF[6][43] ) );
  DFFPOSX1 \RF_reg[6][42]  ( .D(n3837), .CLK(clk), .Q(\RF[6][42] ) );
  DFFPOSX1 \RF_reg[6][41]  ( .D(n3836), .CLK(clk), .Q(\RF[6][41] ) );
  DFFPOSX1 \RF_reg[6][40]  ( .D(n3835), .CLK(clk), .Q(\RF[6][40] ) );
  DFFPOSX1 \RF_reg[6][39]  ( .D(n3834), .CLK(clk), .Q(\RF[6][39] ) );
  DFFPOSX1 \RF_reg[6][38]  ( .D(n3833), .CLK(clk), .Q(\RF[6][38] ) );
  DFFPOSX1 \RF_reg[6][37]  ( .D(n3832), .CLK(clk), .Q(\RF[6][37] ) );
  DFFPOSX1 \RF_reg[6][36]  ( .D(n3831), .CLK(clk), .Q(\RF[6][36] ) );
  DFFPOSX1 \RF_reg[6][35]  ( .D(n3830), .CLK(clk), .Q(\RF[6][35] ) );
  DFFPOSX1 \RF_reg[6][34]  ( .D(n3829), .CLK(clk), .Q(\RF[6][34] ) );
  DFFPOSX1 \RF_reg[6][33]  ( .D(n3828), .CLK(clk), .Q(\RF[6][33] ) );
  DFFPOSX1 \RF_reg[6][32]  ( .D(n3827), .CLK(clk), .Q(\RF[6][32] ) );
  DFFPOSX1 \RF_reg[6][31]  ( .D(n3826), .CLK(clk), .Q(\RF[6][31] ) );
  DFFPOSX1 \RF_reg[6][30]  ( .D(n3825), .CLK(clk), .Q(\RF[6][30] ) );
  DFFPOSX1 \RF_reg[6][29]  ( .D(n3824), .CLK(clk), .Q(\RF[6][29] ) );
  DFFPOSX1 \RF_reg[6][28]  ( .D(n3823), .CLK(clk), .Q(\RF[6][28] ) );
  DFFPOSX1 \RF_reg[6][27]  ( .D(n3822), .CLK(clk), .Q(\RF[6][27] ) );
  DFFPOSX1 \RF_reg[6][26]  ( .D(n3821), .CLK(clk), .Q(\RF[6][26] ) );
  DFFPOSX1 \RF_reg[6][25]  ( .D(n3820), .CLK(clk), .Q(\RF[6][25] ) );
  DFFPOSX1 \RF_reg[6][24]  ( .D(n3819), .CLK(clk), .Q(\RF[6][24] ) );
  DFFPOSX1 \RF_reg[6][23]  ( .D(n3818), .CLK(clk), .Q(\RF[6][23] ) );
  DFFPOSX1 \RF_reg[6][22]  ( .D(n3817), .CLK(clk), .Q(\RF[6][22] ) );
  DFFPOSX1 \RF_reg[6][21]  ( .D(n3816), .CLK(clk), .Q(\RF[6][21] ) );
  DFFPOSX1 \RF_reg[6][20]  ( .D(n3815), .CLK(clk), .Q(\RF[6][20] ) );
  DFFPOSX1 \RF_reg[6][19]  ( .D(n3814), .CLK(clk), .Q(\RF[6][19] ) );
  DFFPOSX1 \RF_reg[6][18]  ( .D(n3813), .CLK(clk), .Q(\RF[6][18] ) );
  DFFPOSX1 \RF_reg[6][17]  ( .D(n3812), .CLK(clk), .Q(\RF[6][17] ) );
  DFFPOSX1 \RF_reg[6][16]  ( .D(n3811), .CLK(clk), .Q(\RF[6][16] ) );
  DFFPOSX1 \RF_reg[6][15]  ( .D(n3810), .CLK(clk), .Q(\RF[6][15] ) );
  DFFPOSX1 \RF_reg[6][14]  ( .D(n3809), .CLK(clk), .Q(\RF[6][14] ) );
  DFFPOSX1 \RF_reg[6][13]  ( .D(n3808), .CLK(clk), .Q(\RF[6][13] ) );
  DFFPOSX1 \RF_reg[6][12]  ( .D(n3807), .CLK(clk), .Q(\RF[6][12] ) );
  DFFPOSX1 \RF_reg[6][11]  ( .D(n3806), .CLK(clk), .Q(\RF[6][11] ) );
  DFFPOSX1 \RF_reg[6][10]  ( .D(n3805), .CLK(clk), .Q(\RF[6][10] ) );
  DFFPOSX1 \RF_reg[6][9]  ( .D(n3804), .CLK(clk), .Q(\RF[6][9] ) );
  DFFPOSX1 \RF_reg[6][8]  ( .D(n3803), .CLK(clk), .Q(\RF[6][8] ) );
  DFFPOSX1 \RF_reg[6][7]  ( .D(n3802), .CLK(clk), .Q(\RF[6][7] ) );
  DFFPOSX1 \RF_reg[6][6]  ( .D(n3801), .CLK(clk), .Q(\RF[6][6] ) );
  DFFPOSX1 \RF_reg[6][5]  ( .D(n3800), .CLK(clk), .Q(\RF[6][5] ) );
  DFFPOSX1 \RF_reg[6][4]  ( .D(n3799), .CLK(clk), .Q(\RF[6][4] ) );
  DFFPOSX1 \RF_reg[6][3]  ( .D(n3798), .CLK(clk), .Q(\RF[6][3] ) );
  DFFPOSX1 \RF_reg[6][2]  ( .D(n3797), .CLK(clk), .Q(\RF[6][2] ) );
  DFFPOSX1 \RF_reg[6][1]  ( .D(n3796), .CLK(clk), .Q(\RF[6][1] ) );
  DFFPOSX1 \RF_reg[6][0]  ( .D(n3795), .CLK(clk), .Q(\RF[6][0] ) );
  DFFPOSX1 \RF_reg[7][63]  ( .D(n3794), .CLK(clk), .Q(\RF[7][63] ) );
  DFFPOSX1 \RF_reg[7][62]  ( .D(n3793), .CLK(clk), .Q(\RF[7][62] ) );
  DFFPOSX1 \RF_reg[7][61]  ( .D(n3792), .CLK(clk), .Q(\RF[7][61] ) );
  DFFPOSX1 \RF_reg[7][60]  ( .D(n3791), .CLK(clk), .Q(\RF[7][60] ) );
  DFFPOSX1 \RF_reg[7][59]  ( .D(n3790), .CLK(clk), .Q(\RF[7][59] ) );
  DFFPOSX1 \RF_reg[7][58]  ( .D(n3789), .CLK(clk), .Q(\RF[7][58] ) );
  DFFPOSX1 \RF_reg[7][57]  ( .D(n3788), .CLK(clk), .Q(\RF[7][57] ) );
  DFFPOSX1 \RF_reg[7][56]  ( .D(n3787), .CLK(clk), .Q(\RF[7][56] ) );
  DFFPOSX1 \RF_reg[7][55]  ( .D(n3786), .CLK(clk), .Q(\RF[7][55] ) );
  DFFPOSX1 \RF_reg[7][54]  ( .D(n3785), .CLK(clk), .Q(\RF[7][54] ) );
  DFFPOSX1 \RF_reg[7][53]  ( .D(n3784), .CLK(clk), .Q(\RF[7][53] ) );
  DFFPOSX1 \RF_reg[7][52]  ( .D(n3783), .CLK(clk), .Q(\RF[7][52] ) );
  DFFPOSX1 \RF_reg[7][51]  ( .D(n3782), .CLK(clk), .Q(\RF[7][51] ) );
  DFFPOSX1 \RF_reg[7][50]  ( .D(n3781), .CLK(clk), .Q(\RF[7][50] ) );
  DFFPOSX1 \RF_reg[7][49]  ( .D(n3780), .CLK(clk), .Q(\RF[7][49] ) );
  DFFPOSX1 \RF_reg[7][48]  ( .D(n3779), .CLK(clk), .Q(\RF[7][48] ) );
  DFFPOSX1 \RF_reg[7][47]  ( .D(n3778), .CLK(clk), .Q(\RF[7][47] ) );
  DFFPOSX1 \RF_reg[7][46]  ( .D(n3777), .CLK(clk), .Q(\RF[7][46] ) );
  DFFPOSX1 \RF_reg[7][45]  ( .D(n3776), .CLK(clk), .Q(\RF[7][45] ) );
  DFFPOSX1 \RF_reg[7][44]  ( .D(n3775), .CLK(clk), .Q(\RF[7][44] ) );
  DFFPOSX1 \RF_reg[7][43]  ( .D(n3774), .CLK(clk), .Q(\RF[7][43] ) );
  DFFPOSX1 \RF_reg[7][42]  ( .D(n3773), .CLK(clk), .Q(\RF[7][42] ) );
  DFFPOSX1 \RF_reg[7][41]  ( .D(n3772), .CLK(clk), .Q(\RF[7][41] ) );
  DFFPOSX1 \RF_reg[7][40]  ( .D(n3771), .CLK(clk), .Q(\RF[7][40] ) );
  DFFPOSX1 \RF_reg[7][39]  ( .D(n3770), .CLK(clk), .Q(\RF[7][39] ) );
  DFFPOSX1 \RF_reg[7][38]  ( .D(n3769), .CLK(clk), .Q(\RF[7][38] ) );
  DFFPOSX1 \RF_reg[7][37]  ( .D(n3768), .CLK(clk), .Q(\RF[7][37] ) );
  DFFPOSX1 \RF_reg[7][36]  ( .D(n3767), .CLK(clk), .Q(\RF[7][36] ) );
  DFFPOSX1 \RF_reg[7][35]  ( .D(n3766), .CLK(clk), .Q(\RF[7][35] ) );
  DFFPOSX1 \RF_reg[7][34]  ( .D(n3765), .CLK(clk), .Q(\RF[7][34] ) );
  DFFPOSX1 \RF_reg[7][33]  ( .D(n3764), .CLK(clk), .Q(\RF[7][33] ) );
  DFFPOSX1 \RF_reg[7][32]  ( .D(n3763), .CLK(clk), .Q(\RF[7][32] ) );
  DFFPOSX1 \RF_reg[7][31]  ( .D(n3762), .CLK(clk), .Q(\RF[7][31] ) );
  DFFPOSX1 \RF_reg[7][30]  ( .D(n3761), .CLK(clk), .Q(\RF[7][30] ) );
  DFFPOSX1 \RF_reg[7][29]  ( .D(n3760), .CLK(clk), .Q(\RF[7][29] ) );
  DFFPOSX1 \RF_reg[7][28]  ( .D(n3759), .CLK(clk), .Q(\RF[7][28] ) );
  DFFPOSX1 \RF_reg[7][27]  ( .D(n3758), .CLK(clk), .Q(\RF[7][27] ) );
  DFFPOSX1 \RF_reg[7][26]  ( .D(n3757), .CLK(clk), .Q(\RF[7][26] ) );
  DFFPOSX1 \RF_reg[7][25]  ( .D(n3756), .CLK(clk), .Q(\RF[7][25] ) );
  DFFPOSX1 \RF_reg[7][24]  ( .D(n3755), .CLK(clk), .Q(\RF[7][24] ) );
  DFFPOSX1 \RF_reg[7][23]  ( .D(n3754), .CLK(clk), .Q(\RF[7][23] ) );
  DFFPOSX1 \RF_reg[7][22]  ( .D(n3753), .CLK(clk), .Q(\RF[7][22] ) );
  DFFPOSX1 \RF_reg[7][21]  ( .D(n3752), .CLK(clk), .Q(\RF[7][21] ) );
  DFFPOSX1 \RF_reg[7][20]  ( .D(n3751), .CLK(clk), .Q(\RF[7][20] ) );
  DFFPOSX1 \RF_reg[7][19]  ( .D(n3750), .CLK(clk), .Q(\RF[7][19] ) );
  DFFPOSX1 \RF_reg[7][18]  ( .D(n3749), .CLK(clk), .Q(\RF[7][18] ) );
  DFFPOSX1 \RF_reg[7][17]  ( .D(n3748), .CLK(clk), .Q(\RF[7][17] ) );
  DFFPOSX1 \RF_reg[7][16]  ( .D(n3747), .CLK(clk), .Q(\RF[7][16] ) );
  DFFPOSX1 \RF_reg[7][15]  ( .D(n3746), .CLK(clk), .Q(\RF[7][15] ) );
  DFFPOSX1 \RF_reg[7][14]  ( .D(n3745), .CLK(clk), .Q(\RF[7][14] ) );
  DFFPOSX1 \RF_reg[7][13]  ( .D(n3744), .CLK(clk), .Q(\RF[7][13] ) );
  DFFPOSX1 \RF_reg[7][12]  ( .D(n3743), .CLK(clk), .Q(\RF[7][12] ) );
  DFFPOSX1 \RF_reg[7][11]  ( .D(n3742), .CLK(clk), .Q(\RF[7][11] ) );
  DFFPOSX1 \RF_reg[7][10]  ( .D(n3741), .CLK(clk), .Q(\RF[7][10] ) );
  DFFPOSX1 \RF_reg[7][9]  ( .D(n3740), .CLK(clk), .Q(\RF[7][9] ) );
  DFFPOSX1 \RF_reg[7][8]  ( .D(n3739), .CLK(clk), .Q(\RF[7][8] ) );
  DFFPOSX1 \RF_reg[7][7]  ( .D(n3738), .CLK(clk), .Q(\RF[7][7] ) );
  DFFPOSX1 \RF_reg[7][6]  ( .D(n3737), .CLK(clk), .Q(\RF[7][6] ) );
  DFFPOSX1 \RF_reg[7][5]  ( .D(n3736), .CLK(clk), .Q(\RF[7][5] ) );
  DFFPOSX1 \RF_reg[7][4]  ( .D(n3735), .CLK(clk), .Q(\RF[7][4] ) );
  DFFPOSX1 \RF_reg[7][3]  ( .D(n3734), .CLK(clk), .Q(\RF[7][3] ) );
  DFFPOSX1 \RF_reg[7][2]  ( .D(n3733), .CLK(clk), .Q(\RF[7][2] ) );
  DFFPOSX1 \RF_reg[7][1]  ( .D(n3732), .CLK(clk), .Q(\RF[7][1] ) );
  DFFPOSX1 \RF_reg[7][0]  ( .D(n3731), .CLK(clk), .Q(\RF[7][0] ) );
  DFFPOSX1 \RF_reg[8][63]  ( .D(n3730), .CLK(clk), .Q(\RF[8][63] ) );
  DFFPOSX1 \RF_reg[8][62]  ( .D(n3729), .CLK(clk), .Q(\RF[8][62] ) );
  DFFPOSX1 \RF_reg[8][61]  ( .D(n3728), .CLK(clk), .Q(\RF[8][61] ) );
  DFFPOSX1 \RF_reg[8][60]  ( .D(n3727), .CLK(clk), .Q(\RF[8][60] ) );
  DFFPOSX1 \RF_reg[8][59]  ( .D(n3726), .CLK(clk), .Q(\RF[8][59] ) );
  DFFPOSX1 \RF_reg[8][58]  ( .D(n3725), .CLK(clk), .Q(\RF[8][58] ) );
  DFFPOSX1 \RF_reg[8][57]  ( .D(n3724), .CLK(clk), .Q(\RF[8][57] ) );
  DFFPOSX1 \RF_reg[8][56]  ( .D(n3723), .CLK(clk), .Q(\RF[8][56] ) );
  DFFPOSX1 \RF_reg[8][55]  ( .D(n3722), .CLK(clk), .Q(\RF[8][55] ) );
  DFFPOSX1 \RF_reg[8][54]  ( .D(n3721), .CLK(clk), .Q(\RF[8][54] ) );
  DFFPOSX1 \RF_reg[8][53]  ( .D(n3720), .CLK(clk), .Q(\RF[8][53] ) );
  DFFPOSX1 \RF_reg[8][52]  ( .D(n3719), .CLK(clk), .Q(\RF[8][52] ) );
  DFFPOSX1 \RF_reg[8][51]  ( .D(n3718), .CLK(clk), .Q(\RF[8][51] ) );
  DFFPOSX1 \RF_reg[8][50]  ( .D(n3717), .CLK(clk), .Q(\RF[8][50] ) );
  DFFPOSX1 \RF_reg[8][49]  ( .D(n3716), .CLK(clk), .Q(\RF[8][49] ) );
  DFFPOSX1 \RF_reg[8][48]  ( .D(n3715), .CLK(clk), .Q(\RF[8][48] ) );
  DFFPOSX1 \RF_reg[8][47]  ( .D(n3714), .CLK(clk), .Q(\RF[8][47] ) );
  DFFPOSX1 \RF_reg[8][46]  ( .D(n3713), .CLK(clk), .Q(\RF[8][46] ) );
  DFFPOSX1 \RF_reg[8][45]  ( .D(n3712), .CLK(clk), .Q(\RF[8][45] ) );
  DFFPOSX1 \RF_reg[8][44]  ( .D(n3711), .CLK(clk), .Q(\RF[8][44] ) );
  DFFPOSX1 \RF_reg[8][43]  ( .D(n3710), .CLK(clk), .Q(\RF[8][43] ) );
  DFFPOSX1 \RF_reg[8][42]  ( .D(n3709), .CLK(clk), .Q(\RF[8][42] ) );
  DFFPOSX1 \RF_reg[8][41]  ( .D(n3708), .CLK(clk), .Q(\RF[8][41] ) );
  DFFPOSX1 \RF_reg[8][40]  ( .D(n3707), .CLK(clk), .Q(\RF[8][40] ) );
  DFFPOSX1 \RF_reg[8][39]  ( .D(n3706), .CLK(clk), .Q(\RF[8][39] ) );
  DFFPOSX1 \RF_reg[8][38]  ( .D(n3705), .CLK(clk), .Q(\RF[8][38] ) );
  DFFPOSX1 \RF_reg[8][37]  ( .D(n3704), .CLK(clk), .Q(\RF[8][37] ) );
  DFFPOSX1 \RF_reg[8][36]  ( .D(n3703), .CLK(clk), .Q(\RF[8][36] ) );
  DFFPOSX1 \RF_reg[8][35]  ( .D(n3702), .CLK(clk), .Q(\RF[8][35] ) );
  DFFPOSX1 \RF_reg[8][34]  ( .D(n3701), .CLK(clk), .Q(\RF[8][34] ) );
  DFFPOSX1 \RF_reg[8][33]  ( .D(n3700), .CLK(clk), .Q(\RF[8][33] ) );
  DFFPOSX1 \RF_reg[8][32]  ( .D(n3699), .CLK(clk), .Q(\RF[8][32] ) );
  DFFPOSX1 \RF_reg[8][31]  ( .D(n3698), .CLK(clk), .Q(\RF[8][31] ) );
  DFFPOSX1 \RF_reg[8][30]  ( .D(n3697), .CLK(clk), .Q(\RF[8][30] ) );
  DFFPOSX1 \RF_reg[8][29]  ( .D(n3696), .CLK(clk), .Q(\RF[8][29] ) );
  DFFPOSX1 \RF_reg[8][28]  ( .D(n3695), .CLK(clk), .Q(\RF[8][28] ) );
  DFFPOSX1 \RF_reg[8][27]  ( .D(n3694), .CLK(clk), .Q(\RF[8][27] ) );
  DFFPOSX1 \RF_reg[8][26]  ( .D(n3693), .CLK(clk), .Q(\RF[8][26] ) );
  DFFPOSX1 \RF_reg[8][25]  ( .D(n3692), .CLK(clk), .Q(\RF[8][25] ) );
  DFFPOSX1 \RF_reg[8][24]  ( .D(n3691), .CLK(clk), .Q(\RF[8][24] ) );
  DFFPOSX1 \RF_reg[8][23]  ( .D(n3690), .CLK(clk), .Q(\RF[8][23] ) );
  DFFPOSX1 \RF_reg[8][22]  ( .D(n3689), .CLK(clk), .Q(\RF[8][22] ) );
  DFFPOSX1 \RF_reg[8][21]  ( .D(n3688), .CLK(clk), .Q(\RF[8][21] ) );
  DFFPOSX1 \RF_reg[8][20]  ( .D(n3687), .CLK(clk), .Q(\RF[8][20] ) );
  DFFPOSX1 \RF_reg[8][19]  ( .D(n3686), .CLK(clk), .Q(\RF[8][19] ) );
  DFFPOSX1 \RF_reg[8][18]  ( .D(n3685), .CLK(clk), .Q(\RF[8][18] ) );
  DFFPOSX1 \RF_reg[8][17]  ( .D(n3684), .CLK(clk), .Q(\RF[8][17] ) );
  DFFPOSX1 \RF_reg[8][16]  ( .D(n3683), .CLK(clk), .Q(\RF[8][16] ) );
  DFFPOSX1 \RF_reg[8][15]  ( .D(n3682), .CLK(clk), .Q(\RF[8][15] ) );
  DFFPOSX1 \RF_reg[8][14]  ( .D(n3681), .CLK(clk), .Q(\RF[8][14] ) );
  DFFPOSX1 \RF_reg[8][13]  ( .D(n3680), .CLK(clk), .Q(\RF[8][13] ) );
  DFFPOSX1 \RF_reg[8][12]  ( .D(n3679), .CLK(clk), .Q(\RF[8][12] ) );
  DFFPOSX1 \RF_reg[8][11]  ( .D(n3678), .CLK(clk), .Q(\RF[8][11] ) );
  DFFPOSX1 \RF_reg[8][10]  ( .D(n3677), .CLK(clk), .Q(\RF[8][10] ) );
  DFFPOSX1 \RF_reg[8][9]  ( .D(n3676), .CLK(clk), .Q(\RF[8][9] ) );
  DFFPOSX1 \RF_reg[8][8]  ( .D(n3675), .CLK(clk), .Q(\RF[8][8] ) );
  DFFPOSX1 \RF_reg[8][7]  ( .D(n3674), .CLK(clk), .Q(\RF[8][7] ) );
  DFFPOSX1 \RF_reg[8][6]  ( .D(n3673), .CLK(clk), .Q(\RF[8][6] ) );
  DFFPOSX1 \RF_reg[8][5]  ( .D(n3672), .CLK(clk), .Q(\RF[8][5] ) );
  DFFPOSX1 \RF_reg[8][4]  ( .D(n3671), .CLK(clk), .Q(\RF[8][4] ) );
  DFFPOSX1 \RF_reg[8][3]  ( .D(n3670), .CLK(clk), .Q(\RF[8][3] ) );
  DFFPOSX1 \RF_reg[8][2]  ( .D(n3669), .CLK(clk), .Q(\RF[8][2] ) );
  DFFPOSX1 \RF_reg[8][1]  ( .D(n3668), .CLK(clk), .Q(\RF[8][1] ) );
  DFFPOSX1 \RF_reg[8][0]  ( .D(n3667), .CLK(clk), .Q(\RF[8][0] ) );
  DFFPOSX1 \RF_reg[9][63]  ( .D(n3666), .CLK(clk), .Q(\RF[9][63] ) );
  DFFPOSX1 \RF_reg[9][62]  ( .D(n3665), .CLK(clk), .Q(\RF[9][62] ) );
  DFFPOSX1 \RF_reg[9][61]  ( .D(n3664), .CLK(clk), .Q(\RF[9][61] ) );
  DFFPOSX1 \RF_reg[9][60]  ( .D(n3663), .CLK(clk), .Q(\RF[9][60] ) );
  DFFPOSX1 \RF_reg[9][59]  ( .D(n3662), .CLK(clk), .Q(\RF[9][59] ) );
  DFFPOSX1 \RF_reg[9][58]  ( .D(n3661), .CLK(clk), .Q(\RF[9][58] ) );
  DFFPOSX1 \RF_reg[9][57]  ( .D(n3660), .CLK(clk), .Q(\RF[9][57] ) );
  DFFPOSX1 \RF_reg[9][56]  ( .D(n3659), .CLK(clk), .Q(\RF[9][56] ) );
  DFFPOSX1 \RF_reg[9][55]  ( .D(n3658), .CLK(clk), .Q(\RF[9][55] ) );
  DFFPOSX1 \RF_reg[9][54]  ( .D(n3657), .CLK(clk), .Q(\RF[9][54] ) );
  DFFPOSX1 \RF_reg[9][53]  ( .D(n3656), .CLK(clk), .Q(\RF[9][53] ) );
  DFFPOSX1 \RF_reg[9][52]  ( .D(n3655), .CLK(clk), .Q(\RF[9][52] ) );
  DFFPOSX1 \RF_reg[9][51]  ( .D(n3654), .CLK(clk), .Q(\RF[9][51] ) );
  DFFPOSX1 \RF_reg[9][50]  ( .D(n3653), .CLK(clk), .Q(\RF[9][50] ) );
  DFFPOSX1 \RF_reg[9][49]  ( .D(n3652), .CLK(clk), .Q(\RF[9][49] ) );
  DFFPOSX1 \RF_reg[9][48]  ( .D(n3651), .CLK(clk), .Q(\RF[9][48] ) );
  DFFPOSX1 \RF_reg[9][47]  ( .D(n3650), .CLK(clk), .Q(\RF[9][47] ) );
  DFFPOSX1 \RF_reg[9][46]  ( .D(n3649), .CLK(clk), .Q(\RF[9][46] ) );
  DFFPOSX1 \RF_reg[9][45]  ( .D(n3648), .CLK(clk), .Q(\RF[9][45] ) );
  DFFPOSX1 \RF_reg[9][44]  ( .D(n3647), .CLK(clk), .Q(\RF[9][44] ) );
  DFFPOSX1 \RF_reg[9][43]  ( .D(n3646), .CLK(clk), .Q(\RF[9][43] ) );
  DFFPOSX1 \RF_reg[9][42]  ( .D(n3645), .CLK(clk), .Q(\RF[9][42] ) );
  DFFPOSX1 \RF_reg[9][41]  ( .D(n3644), .CLK(clk), .Q(\RF[9][41] ) );
  DFFPOSX1 \RF_reg[9][40]  ( .D(n3643), .CLK(clk), .Q(\RF[9][40] ) );
  DFFPOSX1 \RF_reg[9][39]  ( .D(n3642), .CLK(clk), .Q(\RF[9][39] ) );
  DFFPOSX1 \RF_reg[9][38]  ( .D(n3641), .CLK(clk), .Q(\RF[9][38] ) );
  DFFPOSX1 \RF_reg[9][37]  ( .D(n3640), .CLK(clk), .Q(\RF[9][37] ) );
  DFFPOSX1 \RF_reg[9][36]  ( .D(n3639), .CLK(clk), .Q(\RF[9][36] ) );
  DFFPOSX1 \RF_reg[9][35]  ( .D(n3638), .CLK(clk), .Q(\RF[9][35] ) );
  DFFPOSX1 \RF_reg[9][34]  ( .D(n3637), .CLK(clk), .Q(\RF[9][34] ) );
  DFFPOSX1 \RF_reg[9][33]  ( .D(n3636), .CLK(clk), .Q(\RF[9][33] ) );
  DFFPOSX1 \RF_reg[9][32]  ( .D(n3635), .CLK(clk), .Q(\RF[9][32] ) );
  DFFPOSX1 \RF_reg[9][31]  ( .D(n3634), .CLK(clk), .Q(\RF[9][31] ) );
  DFFPOSX1 \RF_reg[9][30]  ( .D(n3633), .CLK(clk), .Q(\RF[9][30] ) );
  DFFPOSX1 \RF_reg[9][29]  ( .D(n3632), .CLK(clk), .Q(\RF[9][29] ) );
  DFFPOSX1 \RF_reg[9][28]  ( .D(n3631), .CLK(clk), .Q(\RF[9][28] ) );
  DFFPOSX1 \RF_reg[9][27]  ( .D(n3630), .CLK(clk), .Q(\RF[9][27] ) );
  DFFPOSX1 \RF_reg[9][26]  ( .D(n3629), .CLK(clk), .Q(\RF[9][26] ) );
  DFFPOSX1 \RF_reg[9][25]  ( .D(n3628), .CLK(clk), .Q(\RF[9][25] ) );
  DFFPOSX1 \RF_reg[9][24]  ( .D(n3627), .CLK(clk), .Q(\RF[9][24] ) );
  DFFPOSX1 \RF_reg[9][23]  ( .D(n3626), .CLK(clk), .Q(\RF[9][23] ) );
  DFFPOSX1 \RF_reg[9][22]  ( .D(n3625), .CLK(clk), .Q(\RF[9][22] ) );
  DFFPOSX1 \RF_reg[9][21]  ( .D(n3624), .CLK(clk), .Q(\RF[9][21] ) );
  DFFPOSX1 \RF_reg[9][20]  ( .D(n3623), .CLK(clk), .Q(\RF[9][20] ) );
  DFFPOSX1 \RF_reg[9][19]  ( .D(n3622), .CLK(clk), .Q(\RF[9][19] ) );
  DFFPOSX1 \RF_reg[9][18]  ( .D(n3621), .CLK(clk), .Q(\RF[9][18] ) );
  DFFPOSX1 \RF_reg[9][17]  ( .D(n3620), .CLK(clk), .Q(\RF[9][17] ) );
  DFFPOSX1 \RF_reg[9][16]  ( .D(n3619), .CLK(clk), .Q(\RF[9][16] ) );
  DFFPOSX1 \RF_reg[9][15]  ( .D(n3618), .CLK(clk), .Q(\RF[9][15] ) );
  DFFPOSX1 \RF_reg[9][14]  ( .D(n3617), .CLK(clk), .Q(\RF[9][14] ) );
  DFFPOSX1 \RF_reg[9][13]  ( .D(n3616), .CLK(clk), .Q(\RF[9][13] ) );
  DFFPOSX1 \RF_reg[9][12]  ( .D(n3615), .CLK(clk), .Q(\RF[9][12] ) );
  DFFPOSX1 \RF_reg[9][11]  ( .D(n3614), .CLK(clk), .Q(\RF[9][11] ) );
  DFFPOSX1 \RF_reg[9][10]  ( .D(n3613), .CLK(clk), .Q(\RF[9][10] ) );
  DFFPOSX1 \RF_reg[9][9]  ( .D(n3612), .CLK(clk), .Q(\RF[9][9] ) );
  DFFPOSX1 \RF_reg[9][8]  ( .D(n3611), .CLK(clk), .Q(\RF[9][8] ) );
  DFFPOSX1 \RF_reg[9][7]  ( .D(n3610), .CLK(clk), .Q(\RF[9][7] ) );
  DFFPOSX1 \RF_reg[9][6]  ( .D(n3609), .CLK(clk), .Q(\RF[9][6] ) );
  DFFPOSX1 \RF_reg[9][5]  ( .D(n3608), .CLK(clk), .Q(\RF[9][5] ) );
  DFFPOSX1 \RF_reg[9][4]  ( .D(n3607), .CLK(clk), .Q(\RF[9][4] ) );
  DFFPOSX1 \RF_reg[9][3]  ( .D(n3606), .CLK(clk), .Q(\RF[9][3] ) );
  DFFPOSX1 \RF_reg[9][2]  ( .D(n3605), .CLK(clk), .Q(\RF[9][2] ) );
  DFFPOSX1 \RF_reg[9][1]  ( .D(n3604), .CLK(clk), .Q(\RF[9][1] ) );
  DFFPOSX1 \RF_reg[9][0]  ( .D(n3603), .CLK(clk), .Q(\RF[9][0] ) );
  DFFPOSX1 \RF_reg[10][63]  ( .D(n3602), .CLK(clk), .Q(\RF[10][63] ) );
  DFFPOSX1 \RF_reg[10][62]  ( .D(n3601), .CLK(clk), .Q(\RF[10][62] ) );
  DFFPOSX1 \RF_reg[10][61]  ( .D(n3600), .CLK(clk), .Q(\RF[10][61] ) );
  DFFPOSX1 \RF_reg[10][60]  ( .D(n3599), .CLK(clk), .Q(\RF[10][60] ) );
  DFFPOSX1 \RF_reg[10][59]  ( .D(n3598), .CLK(clk), .Q(\RF[10][59] ) );
  DFFPOSX1 \RF_reg[10][58]  ( .D(n3597), .CLK(clk), .Q(\RF[10][58] ) );
  DFFPOSX1 \RF_reg[10][57]  ( .D(n3596), .CLK(clk), .Q(\RF[10][57] ) );
  DFFPOSX1 \RF_reg[10][56]  ( .D(n3595), .CLK(clk), .Q(\RF[10][56] ) );
  DFFPOSX1 \RF_reg[10][55]  ( .D(n3594), .CLK(clk), .Q(\RF[10][55] ) );
  DFFPOSX1 \RF_reg[10][54]  ( .D(n3593), .CLK(clk), .Q(\RF[10][54] ) );
  DFFPOSX1 \RF_reg[10][53]  ( .D(n3592), .CLK(clk), .Q(\RF[10][53] ) );
  DFFPOSX1 \RF_reg[10][52]  ( .D(n3591), .CLK(clk), .Q(\RF[10][52] ) );
  DFFPOSX1 \RF_reg[10][51]  ( .D(n3590), .CLK(clk), .Q(\RF[10][51] ) );
  DFFPOSX1 \RF_reg[10][50]  ( .D(n3589), .CLK(clk), .Q(\RF[10][50] ) );
  DFFPOSX1 \RF_reg[10][49]  ( .D(n3588), .CLK(clk), .Q(\RF[10][49] ) );
  DFFPOSX1 \RF_reg[10][48]  ( .D(n3587), .CLK(clk), .Q(\RF[10][48] ) );
  DFFPOSX1 \RF_reg[10][47]  ( .D(n3586), .CLK(clk), .Q(\RF[10][47] ) );
  DFFPOSX1 \RF_reg[10][46]  ( .D(n3585), .CLK(clk), .Q(\RF[10][46] ) );
  DFFPOSX1 \RF_reg[10][45]  ( .D(n3584), .CLK(clk), .Q(\RF[10][45] ) );
  DFFPOSX1 \RF_reg[10][44]  ( .D(n3583), .CLK(clk), .Q(\RF[10][44] ) );
  DFFPOSX1 \RF_reg[10][43]  ( .D(n3582), .CLK(clk), .Q(\RF[10][43] ) );
  DFFPOSX1 \RF_reg[10][42]  ( .D(n3581), .CLK(clk), .Q(\RF[10][42] ) );
  DFFPOSX1 \RF_reg[10][41]  ( .D(n3580), .CLK(clk), .Q(\RF[10][41] ) );
  DFFPOSX1 \RF_reg[10][40]  ( .D(n3579), .CLK(clk), .Q(\RF[10][40] ) );
  DFFPOSX1 \RF_reg[10][39]  ( .D(n3578), .CLK(clk), .Q(\RF[10][39] ) );
  DFFPOSX1 \RF_reg[10][38]  ( .D(n3577), .CLK(clk), .Q(\RF[10][38] ) );
  DFFPOSX1 \RF_reg[10][37]  ( .D(n3576), .CLK(clk), .Q(\RF[10][37] ) );
  DFFPOSX1 \RF_reg[10][36]  ( .D(n3575), .CLK(clk), .Q(\RF[10][36] ) );
  DFFPOSX1 \RF_reg[10][35]  ( .D(n3574), .CLK(clk), .Q(\RF[10][35] ) );
  DFFPOSX1 \RF_reg[10][34]  ( .D(n3573), .CLK(clk), .Q(\RF[10][34] ) );
  DFFPOSX1 \RF_reg[10][33]  ( .D(n3572), .CLK(clk), .Q(\RF[10][33] ) );
  DFFPOSX1 \RF_reg[10][32]  ( .D(n3571), .CLK(clk), .Q(\RF[10][32] ) );
  DFFPOSX1 \RF_reg[10][31]  ( .D(n3570), .CLK(clk), .Q(\RF[10][31] ) );
  DFFPOSX1 \RF_reg[10][30]  ( .D(n3569), .CLK(clk), .Q(\RF[10][30] ) );
  DFFPOSX1 \RF_reg[10][29]  ( .D(n3568), .CLK(clk), .Q(\RF[10][29] ) );
  DFFPOSX1 \RF_reg[10][28]  ( .D(n3567), .CLK(clk), .Q(\RF[10][28] ) );
  DFFPOSX1 \RF_reg[10][27]  ( .D(n3566), .CLK(clk), .Q(\RF[10][27] ) );
  DFFPOSX1 \RF_reg[10][26]  ( .D(n3565), .CLK(clk), .Q(\RF[10][26] ) );
  DFFPOSX1 \RF_reg[10][25]  ( .D(n3564), .CLK(clk), .Q(\RF[10][25] ) );
  DFFPOSX1 \RF_reg[10][24]  ( .D(n3563), .CLK(clk), .Q(\RF[10][24] ) );
  DFFPOSX1 \RF_reg[10][23]  ( .D(n3562), .CLK(clk), .Q(\RF[10][23] ) );
  DFFPOSX1 \RF_reg[10][22]  ( .D(n3561), .CLK(clk), .Q(\RF[10][22] ) );
  DFFPOSX1 \RF_reg[10][21]  ( .D(n3560), .CLK(clk), .Q(\RF[10][21] ) );
  DFFPOSX1 \RF_reg[10][20]  ( .D(n3559), .CLK(clk), .Q(\RF[10][20] ) );
  DFFPOSX1 \RF_reg[10][19]  ( .D(n3558), .CLK(clk), .Q(\RF[10][19] ) );
  DFFPOSX1 \RF_reg[10][18]  ( .D(n3557), .CLK(clk), .Q(\RF[10][18] ) );
  DFFPOSX1 \RF_reg[10][17]  ( .D(n3556), .CLK(clk), .Q(\RF[10][17] ) );
  DFFPOSX1 \RF_reg[10][16]  ( .D(n3555), .CLK(clk), .Q(\RF[10][16] ) );
  DFFPOSX1 \RF_reg[10][15]  ( .D(n3554), .CLK(clk), .Q(\RF[10][15] ) );
  DFFPOSX1 \RF_reg[10][14]  ( .D(n3553), .CLK(clk), .Q(\RF[10][14] ) );
  DFFPOSX1 \RF_reg[10][13]  ( .D(n3552), .CLK(clk), .Q(\RF[10][13] ) );
  DFFPOSX1 \RF_reg[10][12]  ( .D(n3551), .CLK(clk), .Q(\RF[10][12] ) );
  DFFPOSX1 \RF_reg[10][11]  ( .D(n3550), .CLK(clk), .Q(\RF[10][11] ) );
  DFFPOSX1 \RF_reg[10][10]  ( .D(n3549), .CLK(clk), .Q(\RF[10][10] ) );
  DFFPOSX1 \RF_reg[10][9]  ( .D(n3548), .CLK(clk), .Q(\RF[10][9] ) );
  DFFPOSX1 \RF_reg[10][8]  ( .D(n3547), .CLK(clk), .Q(\RF[10][8] ) );
  DFFPOSX1 \RF_reg[10][7]  ( .D(n3546), .CLK(clk), .Q(\RF[10][7] ) );
  DFFPOSX1 \RF_reg[10][6]  ( .D(n3545), .CLK(clk), .Q(\RF[10][6] ) );
  DFFPOSX1 \RF_reg[10][5]  ( .D(n3544), .CLK(clk), .Q(\RF[10][5] ) );
  DFFPOSX1 \RF_reg[10][4]  ( .D(n3543), .CLK(clk), .Q(\RF[10][4] ) );
  DFFPOSX1 \RF_reg[10][3]  ( .D(n3542), .CLK(clk), .Q(\RF[10][3] ) );
  DFFPOSX1 \RF_reg[10][2]  ( .D(n3541), .CLK(clk), .Q(\RF[10][2] ) );
  DFFPOSX1 \RF_reg[10][1]  ( .D(n3540), .CLK(clk), .Q(\RF[10][1] ) );
  DFFPOSX1 \RF_reg[10][0]  ( .D(n3539), .CLK(clk), .Q(\RF[10][0] ) );
  DFFPOSX1 \RF_reg[11][63]  ( .D(n3538), .CLK(clk), .Q(\RF[11][63] ) );
  DFFPOSX1 \RF_reg[11][62]  ( .D(n3537), .CLK(clk), .Q(\RF[11][62] ) );
  DFFPOSX1 \RF_reg[11][61]  ( .D(n3536), .CLK(clk), .Q(\RF[11][61] ) );
  DFFPOSX1 \RF_reg[11][60]  ( .D(n3535), .CLK(clk), .Q(\RF[11][60] ) );
  DFFPOSX1 \RF_reg[11][59]  ( .D(n3534), .CLK(clk), .Q(\RF[11][59] ) );
  DFFPOSX1 \RF_reg[11][58]  ( .D(n3533), .CLK(clk), .Q(\RF[11][58] ) );
  DFFPOSX1 \RF_reg[11][57]  ( .D(n3532), .CLK(clk), .Q(\RF[11][57] ) );
  DFFPOSX1 \RF_reg[11][56]  ( .D(n3531), .CLK(clk), .Q(\RF[11][56] ) );
  DFFPOSX1 \RF_reg[11][55]  ( .D(n3530), .CLK(clk), .Q(\RF[11][55] ) );
  DFFPOSX1 \RF_reg[11][54]  ( .D(n3529), .CLK(clk), .Q(\RF[11][54] ) );
  DFFPOSX1 \RF_reg[11][53]  ( .D(n3528), .CLK(clk), .Q(\RF[11][53] ) );
  DFFPOSX1 \RF_reg[11][52]  ( .D(n3527), .CLK(clk), .Q(\RF[11][52] ) );
  DFFPOSX1 \RF_reg[11][51]  ( .D(n3526), .CLK(clk), .Q(\RF[11][51] ) );
  DFFPOSX1 \RF_reg[11][50]  ( .D(n3525), .CLK(clk), .Q(\RF[11][50] ) );
  DFFPOSX1 \RF_reg[11][49]  ( .D(n3524), .CLK(clk), .Q(\RF[11][49] ) );
  DFFPOSX1 \RF_reg[11][48]  ( .D(n3523), .CLK(clk), .Q(\RF[11][48] ) );
  DFFPOSX1 \RF_reg[11][47]  ( .D(n3522), .CLK(clk), .Q(\RF[11][47] ) );
  DFFPOSX1 \RF_reg[11][46]  ( .D(n3521), .CLK(clk), .Q(\RF[11][46] ) );
  DFFPOSX1 \RF_reg[11][45]  ( .D(n3520), .CLK(clk), .Q(\RF[11][45] ) );
  DFFPOSX1 \RF_reg[11][44]  ( .D(n3519), .CLK(clk), .Q(\RF[11][44] ) );
  DFFPOSX1 \RF_reg[11][43]  ( .D(n3518), .CLK(clk), .Q(\RF[11][43] ) );
  DFFPOSX1 \RF_reg[11][42]  ( .D(n3517), .CLK(clk), .Q(\RF[11][42] ) );
  DFFPOSX1 \RF_reg[11][41]  ( .D(n3516), .CLK(clk), .Q(\RF[11][41] ) );
  DFFPOSX1 \RF_reg[11][40]  ( .D(n3515), .CLK(clk), .Q(\RF[11][40] ) );
  DFFPOSX1 \RF_reg[11][39]  ( .D(n3514), .CLK(clk), .Q(\RF[11][39] ) );
  DFFPOSX1 \RF_reg[11][38]  ( .D(n3513), .CLK(clk), .Q(\RF[11][38] ) );
  DFFPOSX1 \RF_reg[11][37]  ( .D(n3512), .CLK(clk), .Q(\RF[11][37] ) );
  DFFPOSX1 \RF_reg[11][36]  ( .D(n3511), .CLK(clk), .Q(\RF[11][36] ) );
  DFFPOSX1 \RF_reg[11][35]  ( .D(n3510), .CLK(clk), .Q(\RF[11][35] ) );
  DFFPOSX1 \RF_reg[11][34]  ( .D(n3509), .CLK(clk), .Q(\RF[11][34] ) );
  DFFPOSX1 \RF_reg[11][33]  ( .D(n3508), .CLK(clk), .Q(\RF[11][33] ) );
  DFFPOSX1 \RF_reg[11][32]  ( .D(n3507), .CLK(clk), .Q(\RF[11][32] ) );
  DFFPOSX1 \RF_reg[11][31]  ( .D(n3506), .CLK(clk), .Q(\RF[11][31] ) );
  DFFPOSX1 \RF_reg[11][30]  ( .D(n3505), .CLK(clk), .Q(\RF[11][30] ) );
  DFFPOSX1 \RF_reg[11][29]  ( .D(n3504), .CLK(clk), .Q(\RF[11][29] ) );
  DFFPOSX1 \RF_reg[11][28]  ( .D(n3503), .CLK(clk), .Q(\RF[11][28] ) );
  DFFPOSX1 \RF_reg[11][27]  ( .D(n3502), .CLK(clk), .Q(\RF[11][27] ) );
  DFFPOSX1 \RF_reg[11][26]  ( .D(n3501), .CLK(clk), .Q(\RF[11][26] ) );
  DFFPOSX1 \RF_reg[11][25]  ( .D(n3500), .CLK(clk), .Q(\RF[11][25] ) );
  DFFPOSX1 \RF_reg[11][24]  ( .D(n3499), .CLK(clk), .Q(\RF[11][24] ) );
  DFFPOSX1 \RF_reg[11][23]  ( .D(n3498), .CLK(clk), .Q(\RF[11][23] ) );
  DFFPOSX1 \RF_reg[11][22]  ( .D(n3497), .CLK(clk), .Q(\RF[11][22] ) );
  DFFPOSX1 \RF_reg[11][21]  ( .D(n3496), .CLK(clk), .Q(\RF[11][21] ) );
  DFFPOSX1 \RF_reg[11][20]  ( .D(n3495), .CLK(clk), .Q(\RF[11][20] ) );
  DFFPOSX1 \RF_reg[11][19]  ( .D(n3494), .CLK(clk), .Q(\RF[11][19] ) );
  DFFPOSX1 \RF_reg[11][18]  ( .D(n3493), .CLK(clk), .Q(\RF[11][18] ) );
  DFFPOSX1 \RF_reg[11][17]  ( .D(n3492), .CLK(clk), .Q(\RF[11][17] ) );
  DFFPOSX1 \RF_reg[11][16]  ( .D(n3491), .CLK(clk), .Q(\RF[11][16] ) );
  DFFPOSX1 \RF_reg[11][15]  ( .D(n3490), .CLK(clk), .Q(\RF[11][15] ) );
  DFFPOSX1 \RF_reg[11][14]  ( .D(n3489), .CLK(clk), .Q(\RF[11][14] ) );
  DFFPOSX1 \RF_reg[11][13]  ( .D(n3488), .CLK(clk), .Q(\RF[11][13] ) );
  DFFPOSX1 \RF_reg[11][12]  ( .D(n3487), .CLK(clk), .Q(\RF[11][12] ) );
  DFFPOSX1 \RF_reg[11][11]  ( .D(n3486), .CLK(clk), .Q(\RF[11][11] ) );
  DFFPOSX1 \RF_reg[11][10]  ( .D(n3485), .CLK(clk), .Q(\RF[11][10] ) );
  DFFPOSX1 \RF_reg[11][9]  ( .D(n3484), .CLK(clk), .Q(\RF[11][9] ) );
  DFFPOSX1 \RF_reg[11][8]  ( .D(n3483), .CLK(clk), .Q(\RF[11][8] ) );
  DFFPOSX1 \RF_reg[11][7]  ( .D(n3482), .CLK(clk), .Q(\RF[11][7] ) );
  DFFPOSX1 \RF_reg[11][6]  ( .D(n3481), .CLK(clk), .Q(\RF[11][6] ) );
  DFFPOSX1 \RF_reg[11][5]  ( .D(n3480), .CLK(clk), .Q(\RF[11][5] ) );
  DFFPOSX1 \RF_reg[11][4]  ( .D(n3479), .CLK(clk), .Q(\RF[11][4] ) );
  DFFPOSX1 \RF_reg[11][3]  ( .D(n3478), .CLK(clk), .Q(\RF[11][3] ) );
  DFFPOSX1 \RF_reg[11][2]  ( .D(n3477), .CLK(clk), .Q(\RF[11][2] ) );
  DFFPOSX1 \RF_reg[11][1]  ( .D(n3476), .CLK(clk), .Q(\RF[11][1] ) );
  DFFPOSX1 \RF_reg[11][0]  ( .D(n3475), .CLK(clk), .Q(\RF[11][0] ) );
  DFFPOSX1 \RF_reg[12][63]  ( .D(n3474), .CLK(clk), .Q(\RF[12][63] ) );
  DFFPOSX1 \RF_reg[12][62]  ( .D(n3473), .CLK(clk), .Q(\RF[12][62] ) );
  DFFPOSX1 \RF_reg[12][61]  ( .D(n3472), .CLK(clk), .Q(\RF[12][61] ) );
  DFFPOSX1 \RF_reg[12][60]  ( .D(n3471), .CLK(clk), .Q(\RF[12][60] ) );
  DFFPOSX1 \RF_reg[12][59]  ( .D(n3470), .CLK(clk), .Q(\RF[12][59] ) );
  DFFPOSX1 \RF_reg[12][58]  ( .D(n3469), .CLK(clk), .Q(\RF[12][58] ) );
  DFFPOSX1 \RF_reg[12][57]  ( .D(n3468), .CLK(clk), .Q(\RF[12][57] ) );
  DFFPOSX1 \RF_reg[12][56]  ( .D(n3467), .CLK(clk), .Q(\RF[12][56] ) );
  DFFPOSX1 \RF_reg[12][55]  ( .D(n3466), .CLK(clk), .Q(\RF[12][55] ) );
  DFFPOSX1 \RF_reg[12][54]  ( .D(n3465), .CLK(clk), .Q(\RF[12][54] ) );
  DFFPOSX1 \RF_reg[12][53]  ( .D(n3464), .CLK(clk), .Q(\RF[12][53] ) );
  DFFPOSX1 \RF_reg[12][52]  ( .D(n3463), .CLK(clk), .Q(\RF[12][52] ) );
  DFFPOSX1 \RF_reg[12][51]  ( .D(n3462), .CLK(clk), .Q(\RF[12][51] ) );
  DFFPOSX1 \RF_reg[12][50]  ( .D(n3461), .CLK(clk), .Q(\RF[12][50] ) );
  DFFPOSX1 \RF_reg[12][49]  ( .D(n3460), .CLK(clk), .Q(\RF[12][49] ) );
  DFFPOSX1 \RF_reg[12][48]  ( .D(n3459), .CLK(clk), .Q(\RF[12][48] ) );
  DFFPOSX1 \RF_reg[12][47]  ( .D(n3458), .CLK(clk), .Q(\RF[12][47] ) );
  DFFPOSX1 \RF_reg[12][46]  ( .D(n3457), .CLK(clk), .Q(\RF[12][46] ) );
  DFFPOSX1 \RF_reg[12][45]  ( .D(n3456), .CLK(clk), .Q(\RF[12][45] ) );
  DFFPOSX1 \RF_reg[12][44]  ( .D(n3455), .CLK(clk), .Q(\RF[12][44] ) );
  DFFPOSX1 \RF_reg[12][43]  ( .D(n3454), .CLK(clk), .Q(\RF[12][43] ) );
  DFFPOSX1 \RF_reg[12][42]  ( .D(n3453), .CLK(clk), .Q(\RF[12][42] ) );
  DFFPOSX1 \RF_reg[12][41]  ( .D(n3452), .CLK(clk), .Q(\RF[12][41] ) );
  DFFPOSX1 \RF_reg[12][40]  ( .D(n3451), .CLK(clk), .Q(\RF[12][40] ) );
  DFFPOSX1 \RF_reg[12][39]  ( .D(n3450), .CLK(clk), .Q(\RF[12][39] ) );
  DFFPOSX1 \RF_reg[12][38]  ( .D(n3449), .CLK(clk), .Q(\RF[12][38] ) );
  DFFPOSX1 \RF_reg[12][37]  ( .D(n3448), .CLK(clk), .Q(\RF[12][37] ) );
  DFFPOSX1 \RF_reg[12][36]  ( .D(n3447), .CLK(clk), .Q(\RF[12][36] ) );
  DFFPOSX1 \RF_reg[12][35]  ( .D(n3446), .CLK(clk), .Q(\RF[12][35] ) );
  DFFPOSX1 \RF_reg[12][34]  ( .D(n3445), .CLK(clk), .Q(\RF[12][34] ) );
  DFFPOSX1 \RF_reg[12][33]  ( .D(n3444), .CLK(clk), .Q(\RF[12][33] ) );
  DFFPOSX1 \RF_reg[12][32]  ( .D(n3443), .CLK(clk), .Q(\RF[12][32] ) );
  DFFPOSX1 \RF_reg[12][31]  ( .D(n3442), .CLK(clk), .Q(\RF[12][31] ) );
  DFFPOSX1 \RF_reg[12][30]  ( .D(n3441), .CLK(clk), .Q(\RF[12][30] ) );
  DFFPOSX1 \RF_reg[12][29]  ( .D(n3440), .CLK(clk), .Q(\RF[12][29] ) );
  DFFPOSX1 \RF_reg[12][28]  ( .D(n3439), .CLK(clk), .Q(\RF[12][28] ) );
  DFFPOSX1 \RF_reg[12][27]  ( .D(n3438), .CLK(clk), .Q(\RF[12][27] ) );
  DFFPOSX1 \RF_reg[12][26]  ( .D(n3437), .CLK(clk), .Q(\RF[12][26] ) );
  DFFPOSX1 \RF_reg[12][25]  ( .D(n3436), .CLK(clk), .Q(\RF[12][25] ) );
  DFFPOSX1 \RF_reg[12][24]  ( .D(n3435), .CLK(clk), .Q(\RF[12][24] ) );
  DFFPOSX1 \RF_reg[12][23]  ( .D(n3434), .CLK(clk), .Q(\RF[12][23] ) );
  DFFPOSX1 \RF_reg[12][22]  ( .D(n3433), .CLK(clk), .Q(\RF[12][22] ) );
  DFFPOSX1 \RF_reg[12][21]  ( .D(n3432), .CLK(clk), .Q(\RF[12][21] ) );
  DFFPOSX1 \RF_reg[12][20]  ( .D(n3431), .CLK(clk), .Q(\RF[12][20] ) );
  DFFPOSX1 \RF_reg[12][19]  ( .D(n3430), .CLK(clk), .Q(\RF[12][19] ) );
  DFFPOSX1 \RF_reg[12][18]  ( .D(n3429), .CLK(clk), .Q(\RF[12][18] ) );
  DFFPOSX1 \RF_reg[12][17]  ( .D(n3428), .CLK(clk), .Q(\RF[12][17] ) );
  DFFPOSX1 \RF_reg[12][16]  ( .D(n3427), .CLK(clk), .Q(\RF[12][16] ) );
  DFFPOSX1 \RF_reg[12][15]  ( .D(n3426), .CLK(clk), .Q(\RF[12][15] ) );
  DFFPOSX1 \RF_reg[12][14]  ( .D(n3425), .CLK(clk), .Q(\RF[12][14] ) );
  DFFPOSX1 \RF_reg[12][13]  ( .D(n3424), .CLK(clk), .Q(\RF[12][13] ) );
  DFFPOSX1 \RF_reg[12][12]  ( .D(n3423), .CLK(clk), .Q(\RF[12][12] ) );
  DFFPOSX1 \RF_reg[12][11]  ( .D(n3422), .CLK(clk), .Q(\RF[12][11] ) );
  DFFPOSX1 \RF_reg[12][10]  ( .D(n3421), .CLK(clk), .Q(\RF[12][10] ) );
  DFFPOSX1 \RF_reg[12][9]  ( .D(n3420), .CLK(clk), .Q(\RF[12][9] ) );
  DFFPOSX1 \RF_reg[12][8]  ( .D(n3419), .CLK(clk), .Q(\RF[12][8] ) );
  DFFPOSX1 \RF_reg[12][7]  ( .D(n3418), .CLK(clk), .Q(\RF[12][7] ) );
  DFFPOSX1 \RF_reg[12][6]  ( .D(n3417), .CLK(clk), .Q(\RF[12][6] ) );
  DFFPOSX1 \RF_reg[12][5]  ( .D(n3416), .CLK(clk), .Q(\RF[12][5] ) );
  DFFPOSX1 \RF_reg[12][4]  ( .D(n3415), .CLK(clk), .Q(\RF[12][4] ) );
  DFFPOSX1 \RF_reg[12][3]  ( .D(n3414), .CLK(clk), .Q(\RF[12][3] ) );
  DFFPOSX1 \RF_reg[12][2]  ( .D(n3413), .CLK(clk), .Q(\RF[12][2] ) );
  DFFPOSX1 \RF_reg[12][1]  ( .D(n3412), .CLK(clk), .Q(\RF[12][1] ) );
  DFFPOSX1 \RF_reg[12][0]  ( .D(n3411), .CLK(clk), .Q(\RF[12][0] ) );
  DFFPOSX1 \RF_reg[13][63]  ( .D(n3410), .CLK(clk), .Q(\RF[13][63] ) );
  DFFPOSX1 \RF_reg[13][62]  ( .D(n3409), .CLK(clk), .Q(\RF[13][62] ) );
  DFFPOSX1 \RF_reg[13][61]  ( .D(n3408), .CLK(clk), .Q(\RF[13][61] ) );
  DFFPOSX1 \RF_reg[13][60]  ( .D(n3407), .CLK(clk), .Q(\RF[13][60] ) );
  DFFPOSX1 \RF_reg[13][59]  ( .D(n3406), .CLK(clk), .Q(\RF[13][59] ) );
  DFFPOSX1 \RF_reg[13][58]  ( .D(n3405), .CLK(clk), .Q(\RF[13][58] ) );
  DFFPOSX1 \RF_reg[13][57]  ( .D(n3404), .CLK(clk), .Q(\RF[13][57] ) );
  DFFPOSX1 \RF_reg[13][56]  ( .D(n3403), .CLK(clk), .Q(\RF[13][56] ) );
  DFFPOSX1 \RF_reg[13][55]  ( .D(n3402), .CLK(clk), .Q(\RF[13][55] ) );
  DFFPOSX1 \RF_reg[13][54]  ( .D(n3401), .CLK(clk), .Q(\RF[13][54] ) );
  DFFPOSX1 \RF_reg[13][53]  ( .D(n3400), .CLK(clk), .Q(\RF[13][53] ) );
  DFFPOSX1 \RF_reg[13][52]  ( .D(n3399), .CLK(clk), .Q(\RF[13][52] ) );
  DFFPOSX1 \RF_reg[13][51]  ( .D(n3398), .CLK(clk), .Q(\RF[13][51] ) );
  DFFPOSX1 \RF_reg[13][50]  ( .D(n3397), .CLK(clk), .Q(\RF[13][50] ) );
  DFFPOSX1 \RF_reg[13][49]  ( .D(n3396), .CLK(clk), .Q(\RF[13][49] ) );
  DFFPOSX1 \RF_reg[13][48]  ( .D(n3395), .CLK(clk), .Q(\RF[13][48] ) );
  DFFPOSX1 \RF_reg[13][47]  ( .D(n3394), .CLK(clk), .Q(\RF[13][47] ) );
  DFFPOSX1 \RF_reg[13][46]  ( .D(n3393), .CLK(clk), .Q(\RF[13][46] ) );
  DFFPOSX1 \RF_reg[13][45]  ( .D(n3392), .CLK(clk), .Q(\RF[13][45] ) );
  DFFPOSX1 \RF_reg[13][44]  ( .D(n3391), .CLK(clk), .Q(\RF[13][44] ) );
  DFFPOSX1 \RF_reg[13][43]  ( .D(n3390), .CLK(clk), .Q(\RF[13][43] ) );
  DFFPOSX1 \RF_reg[13][42]  ( .D(n3389), .CLK(clk), .Q(\RF[13][42] ) );
  DFFPOSX1 \RF_reg[13][41]  ( .D(n3388), .CLK(clk), .Q(\RF[13][41] ) );
  DFFPOSX1 \RF_reg[13][40]  ( .D(n3387), .CLK(clk), .Q(\RF[13][40] ) );
  DFFPOSX1 \RF_reg[13][39]  ( .D(n3386), .CLK(clk), .Q(\RF[13][39] ) );
  DFFPOSX1 \RF_reg[13][38]  ( .D(n3385), .CLK(clk), .Q(\RF[13][38] ) );
  DFFPOSX1 \RF_reg[13][37]  ( .D(n3384), .CLK(clk), .Q(\RF[13][37] ) );
  DFFPOSX1 \RF_reg[13][36]  ( .D(n3383), .CLK(clk), .Q(\RF[13][36] ) );
  DFFPOSX1 \RF_reg[13][35]  ( .D(n3382), .CLK(clk), .Q(\RF[13][35] ) );
  DFFPOSX1 \RF_reg[13][34]  ( .D(n3381), .CLK(clk), .Q(\RF[13][34] ) );
  DFFPOSX1 \RF_reg[13][33]  ( .D(n3380), .CLK(clk), .Q(\RF[13][33] ) );
  DFFPOSX1 \RF_reg[13][32]  ( .D(n3379), .CLK(clk), .Q(\RF[13][32] ) );
  DFFPOSX1 \RF_reg[13][31]  ( .D(n3378), .CLK(clk), .Q(\RF[13][31] ) );
  DFFPOSX1 \RF_reg[13][30]  ( .D(n3377), .CLK(clk), .Q(\RF[13][30] ) );
  DFFPOSX1 \RF_reg[13][29]  ( .D(n3376), .CLK(clk), .Q(\RF[13][29] ) );
  DFFPOSX1 \RF_reg[13][28]  ( .D(n3375), .CLK(clk), .Q(\RF[13][28] ) );
  DFFPOSX1 \RF_reg[13][27]  ( .D(n3374), .CLK(clk), .Q(\RF[13][27] ) );
  DFFPOSX1 \RF_reg[13][26]  ( .D(n3373), .CLK(clk), .Q(\RF[13][26] ) );
  DFFPOSX1 \RF_reg[13][25]  ( .D(n3372), .CLK(clk), .Q(\RF[13][25] ) );
  DFFPOSX1 \RF_reg[13][24]  ( .D(n3371), .CLK(clk), .Q(\RF[13][24] ) );
  DFFPOSX1 \RF_reg[13][23]  ( .D(n3370), .CLK(clk), .Q(\RF[13][23] ) );
  DFFPOSX1 \RF_reg[13][22]  ( .D(n3369), .CLK(clk), .Q(\RF[13][22] ) );
  DFFPOSX1 \RF_reg[13][21]  ( .D(n3368), .CLK(clk), .Q(\RF[13][21] ) );
  DFFPOSX1 \RF_reg[13][20]  ( .D(n3367), .CLK(clk), .Q(\RF[13][20] ) );
  DFFPOSX1 \RF_reg[13][19]  ( .D(n3366), .CLK(clk), .Q(\RF[13][19] ) );
  DFFPOSX1 \RF_reg[13][18]  ( .D(n3365), .CLK(clk), .Q(\RF[13][18] ) );
  DFFPOSX1 \RF_reg[13][17]  ( .D(n3364), .CLK(clk), .Q(\RF[13][17] ) );
  DFFPOSX1 \RF_reg[13][16]  ( .D(n3363), .CLK(clk), .Q(\RF[13][16] ) );
  DFFPOSX1 \RF_reg[13][15]  ( .D(n3362), .CLK(clk), .Q(\RF[13][15] ) );
  DFFPOSX1 \RF_reg[13][14]  ( .D(n3361), .CLK(clk), .Q(\RF[13][14] ) );
  DFFPOSX1 \RF_reg[13][13]  ( .D(n3360), .CLK(clk), .Q(\RF[13][13] ) );
  DFFPOSX1 \RF_reg[13][12]  ( .D(n3359), .CLK(clk), .Q(\RF[13][12] ) );
  DFFPOSX1 \RF_reg[13][11]  ( .D(n3358), .CLK(clk), .Q(\RF[13][11] ) );
  DFFPOSX1 \RF_reg[13][10]  ( .D(n3357), .CLK(clk), .Q(\RF[13][10] ) );
  DFFPOSX1 \RF_reg[13][9]  ( .D(n3356), .CLK(clk), .Q(\RF[13][9] ) );
  DFFPOSX1 \RF_reg[13][8]  ( .D(n3355), .CLK(clk), .Q(\RF[13][8] ) );
  DFFPOSX1 \RF_reg[13][7]  ( .D(n3354), .CLK(clk), .Q(\RF[13][7] ) );
  DFFPOSX1 \RF_reg[13][6]  ( .D(n3353), .CLK(clk), .Q(\RF[13][6] ) );
  DFFPOSX1 \RF_reg[13][5]  ( .D(n3352), .CLK(clk), .Q(\RF[13][5] ) );
  DFFPOSX1 \RF_reg[13][4]  ( .D(n3351), .CLK(clk), .Q(\RF[13][4] ) );
  DFFPOSX1 \RF_reg[13][3]  ( .D(n3350), .CLK(clk), .Q(\RF[13][3] ) );
  DFFPOSX1 \RF_reg[13][2]  ( .D(n3349), .CLK(clk), .Q(\RF[13][2] ) );
  DFFPOSX1 \RF_reg[13][1]  ( .D(n3348), .CLK(clk), .Q(\RF[13][1] ) );
  DFFPOSX1 \RF_reg[13][0]  ( .D(n3347), .CLK(clk), .Q(\RF[13][0] ) );
  DFFPOSX1 \RF_reg[14][63]  ( .D(n3346), .CLK(clk), .Q(\RF[14][63] ) );
  DFFPOSX1 \RF_reg[14][62]  ( .D(n3345), .CLK(clk), .Q(\RF[14][62] ) );
  DFFPOSX1 \RF_reg[14][61]  ( .D(n3344), .CLK(clk), .Q(\RF[14][61] ) );
  DFFPOSX1 \RF_reg[14][60]  ( .D(n3343), .CLK(clk), .Q(\RF[14][60] ) );
  DFFPOSX1 \RF_reg[14][59]  ( .D(n3342), .CLK(clk), .Q(\RF[14][59] ) );
  DFFPOSX1 \RF_reg[14][58]  ( .D(n3341), .CLK(clk), .Q(\RF[14][58] ) );
  DFFPOSX1 \RF_reg[14][57]  ( .D(n3340), .CLK(clk), .Q(\RF[14][57] ) );
  DFFPOSX1 \RF_reg[14][56]  ( .D(n3339), .CLK(clk), .Q(\RF[14][56] ) );
  DFFPOSX1 \RF_reg[14][55]  ( .D(n3338), .CLK(clk), .Q(\RF[14][55] ) );
  DFFPOSX1 \RF_reg[14][54]  ( .D(n3337), .CLK(clk), .Q(\RF[14][54] ) );
  DFFPOSX1 \RF_reg[14][53]  ( .D(n3336), .CLK(clk), .Q(\RF[14][53] ) );
  DFFPOSX1 \RF_reg[14][52]  ( .D(n3335), .CLK(clk), .Q(\RF[14][52] ) );
  DFFPOSX1 \RF_reg[14][51]  ( .D(n3334), .CLK(clk), .Q(\RF[14][51] ) );
  DFFPOSX1 \RF_reg[14][50]  ( .D(n3333), .CLK(clk), .Q(\RF[14][50] ) );
  DFFPOSX1 \RF_reg[14][49]  ( .D(n3332), .CLK(clk), .Q(\RF[14][49] ) );
  DFFPOSX1 \RF_reg[14][48]  ( .D(n3331), .CLK(clk), .Q(\RF[14][48] ) );
  DFFPOSX1 \RF_reg[14][47]  ( .D(n3330), .CLK(clk), .Q(\RF[14][47] ) );
  DFFPOSX1 \RF_reg[14][46]  ( .D(n3329), .CLK(clk), .Q(\RF[14][46] ) );
  DFFPOSX1 \RF_reg[14][45]  ( .D(n3328), .CLK(clk), .Q(\RF[14][45] ) );
  DFFPOSX1 \RF_reg[14][44]  ( .D(n3327), .CLK(clk), .Q(\RF[14][44] ) );
  DFFPOSX1 \RF_reg[14][43]  ( .D(n3326), .CLK(clk), .Q(\RF[14][43] ) );
  DFFPOSX1 \RF_reg[14][42]  ( .D(n3325), .CLK(clk), .Q(\RF[14][42] ) );
  DFFPOSX1 \RF_reg[14][41]  ( .D(n3324), .CLK(clk), .Q(\RF[14][41] ) );
  DFFPOSX1 \RF_reg[14][40]  ( .D(n3323), .CLK(clk), .Q(\RF[14][40] ) );
  DFFPOSX1 \RF_reg[14][39]  ( .D(n3322), .CLK(clk), .Q(\RF[14][39] ) );
  DFFPOSX1 \RF_reg[14][38]  ( .D(n3321), .CLK(clk), .Q(\RF[14][38] ) );
  DFFPOSX1 \RF_reg[14][37]  ( .D(n3320), .CLK(clk), .Q(\RF[14][37] ) );
  DFFPOSX1 \RF_reg[14][36]  ( .D(n3319), .CLK(clk), .Q(\RF[14][36] ) );
  DFFPOSX1 \RF_reg[14][35]  ( .D(n3318), .CLK(clk), .Q(\RF[14][35] ) );
  DFFPOSX1 \RF_reg[14][34]  ( .D(n3317), .CLK(clk), .Q(\RF[14][34] ) );
  DFFPOSX1 \RF_reg[14][33]  ( .D(n3316), .CLK(clk), .Q(\RF[14][33] ) );
  DFFPOSX1 \RF_reg[14][32]  ( .D(n3315), .CLK(clk), .Q(\RF[14][32] ) );
  DFFPOSX1 \RF_reg[14][31]  ( .D(n3314), .CLK(clk), .Q(\RF[14][31] ) );
  DFFPOSX1 \RF_reg[14][30]  ( .D(n3313), .CLK(clk), .Q(\RF[14][30] ) );
  DFFPOSX1 \RF_reg[14][29]  ( .D(n3312), .CLK(clk), .Q(\RF[14][29] ) );
  DFFPOSX1 \RF_reg[14][28]  ( .D(n3311), .CLK(clk), .Q(\RF[14][28] ) );
  DFFPOSX1 \RF_reg[14][27]  ( .D(n3310), .CLK(clk), .Q(\RF[14][27] ) );
  DFFPOSX1 \RF_reg[14][26]  ( .D(n3309), .CLK(clk), .Q(\RF[14][26] ) );
  DFFPOSX1 \RF_reg[14][25]  ( .D(n3308), .CLK(clk), .Q(\RF[14][25] ) );
  DFFPOSX1 \RF_reg[14][24]  ( .D(n3307), .CLK(clk), .Q(\RF[14][24] ) );
  DFFPOSX1 \RF_reg[14][23]  ( .D(n3306), .CLK(clk), .Q(\RF[14][23] ) );
  DFFPOSX1 \RF_reg[14][22]  ( .D(n3305), .CLK(clk), .Q(\RF[14][22] ) );
  DFFPOSX1 \RF_reg[14][21]  ( .D(n3304), .CLK(clk), .Q(\RF[14][21] ) );
  DFFPOSX1 \RF_reg[14][20]  ( .D(n3303), .CLK(clk), .Q(\RF[14][20] ) );
  DFFPOSX1 \RF_reg[14][19]  ( .D(n3302), .CLK(clk), .Q(\RF[14][19] ) );
  DFFPOSX1 \RF_reg[14][18]  ( .D(n3301), .CLK(clk), .Q(\RF[14][18] ) );
  DFFPOSX1 \RF_reg[14][17]  ( .D(n3300), .CLK(clk), .Q(\RF[14][17] ) );
  DFFPOSX1 \RF_reg[14][16]  ( .D(n3299), .CLK(clk), .Q(\RF[14][16] ) );
  DFFPOSX1 \RF_reg[14][15]  ( .D(n3298), .CLK(clk), .Q(\RF[14][15] ) );
  DFFPOSX1 \RF_reg[14][14]  ( .D(n3297), .CLK(clk), .Q(\RF[14][14] ) );
  DFFPOSX1 \RF_reg[14][13]  ( .D(n3296), .CLK(clk), .Q(\RF[14][13] ) );
  DFFPOSX1 \RF_reg[14][12]  ( .D(n3295), .CLK(clk), .Q(\RF[14][12] ) );
  DFFPOSX1 \RF_reg[14][11]  ( .D(n3294), .CLK(clk), .Q(\RF[14][11] ) );
  DFFPOSX1 \RF_reg[14][10]  ( .D(n3293), .CLK(clk), .Q(\RF[14][10] ) );
  DFFPOSX1 \RF_reg[14][9]  ( .D(n3292), .CLK(clk), .Q(\RF[14][9] ) );
  DFFPOSX1 \RF_reg[14][8]  ( .D(n3291), .CLK(clk), .Q(\RF[14][8] ) );
  DFFPOSX1 \RF_reg[14][7]  ( .D(n3290), .CLK(clk), .Q(\RF[14][7] ) );
  DFFPOSX1 \RF_reg[14][6]  ( .D(n3289), .CLK(clk), .Q(\RF[14][6] ) );
  DFFPOSX1 \RF_reg[14][5]  ( .D(n3288), .CLK(clk), .Q(\RF[14][5] ) );
  DFFPOSX1 \RF_reg[14][4]  ( .D(n3287), .CLK(clk), .Q(\RF[14][4] ) );
  DFFPOSX1 \RF_reg[14][3]  ( .D(n3286), .CLK(clk), .Q(\RF[14][3] ) );
  DFFPOSX1 \RF_reg[14][2]  ( .D(n3285), .CLK(clk), .Q(\RF[14][2] ) );
  DFFPOSX1 \RF_reg[14][1]  ( .D(n3284), .CLK(clk), .Q(\RF[14][1] ) );
  DFFPOSX1 \RF_reg[14][0]  ( .D(n3283), .CLK(clk), .Q(\RF[14][0] ) );
  DFFPOSX1 \RF_reg[15][63]  ( .D(n3282), .CLK(clk), .Q(\RF[15][63] ) );
  DFFPOSX1 \RF_reg[15][62]  ( .D(n3281), .CLK(clk), .Q(\RF[15][62] ) );
  DFFPOSX1 \RF_reg[15][61]  ( .D(n3280), .CLK(clk), .Q(\RF[15][61] ) );
  DFFPOSX1 \RF_reg[15][60]  ( .D(n3279), .CLK(clk), .Q(\RF[15][60] ) );
  DFFPOSX1 \RF_reg[15][59]  ( .D(n3278), .CLK(clk), .Q(\RF[15][59] ) );
  DFFPOSX1 \RF_reg[15][58]  ( .D(n3277), .CLK(clk), .Q(\RF[15][58] ) );
  DFFPOSX1 \RF_reg[15][57]  ( .D(n3276), .CLK(clk), .Q(\RF[15][57] ) );
  DFFPOSX1 \RF_reg[15][56]  ( .D(n3275), .CLK(clk), .Q(\RF[15][56] ) );
  DFFPOSX1 \RF_reg[15][55]  ( .D(n3274), .CLK(clk), .Q(\RF[15][55] ) );
  DFFPOSX1 \RF_reg[15][54]  ( .D(n3273), .CLK(clk), .Q(\RF[15][54] ) );
  DFFPOSX1 \RF_reg[15][53]  ( .D(n3272), .CLK(clk), .Q(\RF[15][53] ) );
  DFFPOSX1 \RF_reg[15][52]  ( .D(n3271), .CLK(clk), .Q(\RF[15][52] ) );
  DFFPOSX1 \RF_reg[15][51]  ( .D(n3270), .CLK(clk), .Q(\RF[15][51] ) );
  DFFPOSX1 \RF_reg[15][50]  ( .D(n3269), .CLK(clk), .Q(\RF[15][50] ) );
  DFFPOSX1 \RF_reg[15][49]  ( .D(n3268), .CLK(clk), .Q(\RF[15][49] ) );
  DFFPOSX1 \RF_reg[15][48]  ( .D(n3267), .CLK(clk), .Q(\RF[15][48] ) );
  DFFPOSX1 \RF_reg[15][47]  ( .D(n3266), .CLK(clk), .Q(\RF[15][47] ) );
  DFFPOSX1 \RF_reg[15][46]  ( .D(n3265), .CLK(clk), .Q(\RF[15][46] ) );
  DFFPOSX1 \RF_reg[15][45]  ( .D(n3264), .CLK(clk), .Q(\RF[15][45] ) );
  DFFPOSX1 \RF_reg[15][44]  ( .D(n3263), .CLK(clk), .Q(\RF[15][44] ) );
  DFFPOSX1 \RF_reg[15][43]  ( .D(n3262), .CLK(clk), .Q(\RF[15][43] ) );
  DFFPOSX1 \RF_reg[15][42]  ( .D(n3261), .CLK(clk), .Q(\RF[15][42] ) );
  DFFPOSX1 \RF_reg[15][41]  ( .D(n3260), .CLK(clk), .Q(\RF[15][41] ) );
  DFFPOSX1 \RF_reg[15][40]  ( .D(n3259), .CLK(clk), .Q(\RF[15][40] ) );
  DFFPOSX1 \RF_reg[15][39]  ( .D(n3258), .CLK(clk), .Q(\RF[15][39] ) );
  DFFPOSX1 \RF_reg[15][38]  ( .D(n3257), .CLK(clk), .Q(\RF[15][38] ) );
  DFFPOSX1 \RF_reg[15][37]  ( .D(n3256), .CLK(clk), .Q(\RF[15][37] ) );
  DFFPOSX1 \RF_reg[15][36]  ( .D(n3255), .CLK(clk), .Q(\RF[15][36] ) );
  DFFPOSX1 \RF_reg[15][35]  ( .D(n3254), .CLK(clk), .Q(\RF[15][35] ) );
  DFFPOSX1 \RF_reg[15][34]  ( .D(n3253), .CLK(clk), .Q(\RF[15][34] ) );
  DFFPOSX1 \RF_reg[15][33]  ( .D(n3252), .CLK(clk), .Q(\RF[15][33] ) );
  DFFPOSX1 \RF_reg[15][32]  ( .D(n3251), .CLK(clk), .Q(\RF[15][32] ) );
  DFFPOSX1 \RF_reg[15][31]  ( .D(n3250), .CLK(clk), .Q(\RF[15][31] ) );
  DFFPOSX1 \RF_reg[15][30]  ( .D(n3249), .CLK(clk), .Q(\RF[15][30] ) );
  DFFPOSX1 \RF_reg[15][29]  ( .D(n3248), .CLK(clk), .Q(\RF[15][29] ) );
  DFFPOSX1 \RF_reg[15][28]  ( .D(n3247), .CLK(clk), .Q(\RF[15][28] ) );
  DFFPOSX1 \RF_reg[15][27]  ( .D(n3246), .CLK(clk), .Q(\RF[15][27] ) );
  DFFPOSX1 \RF_reg[15][26]  ( .D(n3245), .CLK(clk), .Q(\RF[15][26] ) );
  DFFPOSX1 \RF_reg[15][25]  ( .D(n3244), .CLK(clk), .Q(\RF[15][25] ) );
  DFFPOSX1 \RF_reg[15][24]  ( .D(n3243), .CLK(clk), .Q(\RF[15][24] ) );
  DFFPOSX1 \RF_reg[15][23]  ( .D(n3242), .CLK(clk), .Q(\RF[15][23] ) );
  DFFPOSX1 \RF_reg[15][22]  ( .D(n3241), .CLK(clk), .Q(\RF[15][22] ) );
  DFFPOSX1 \RF_reg[15][21]  ( .D(n3240), .CLK(clk), .Q(\RF[15][21] ) );
  DFFPOSX1 \RF_reg[15][20]  ( .D(n3239), .CLK(clk), .Q(\RF[15][20] ) );
  DFFPOSX1 \RF_reg[15][19]  ( .D(n3238), .CLK(clk), .Q(\RF[15][19] ) );
  DFFPOSX1 \RF_reg[15][18]  ( .D(n3237), .CLK(clk), .Q(\RF[15][18] ) );
  DFFPOSX1 \RF_reg[15][17]  ( .D(n3236), .CLK(clk), .Q(\RF[15][17] ) );
  DFFPOSX1 \RF_reg[15][16]  ( .D(n3235), .CLK(clk), .Q(\RF[15][16] ) );
  DFFPOSX1 \RF_reg[15][15]  ( .D(n3234), .CLK(clk), .Q(\RF[15][15] ) );
  DFFPOSX1 \RF_reg[15][14]  ( .D(n3233), .CLK(clk), .Q(\RF[15][14] ) );
  DFFPOSX1 \RF_reg[15][13]  ( .D(n3232), .CLK(clk), .Q(\RF[15][13] ) );
  DFFPOSX1 \RF_reg[15][12]  ( .D(n3231), .CLK(clk), .Q(\RF[15][12] ) );
  DFFPOSX1 \RF_reg[15][11]  ( .D(n3230), .CLK(clk), .Q(\RF[15][11] ) );
  DFFPOSX1 \RF_reg[15][10]  ( .D(n3229), .CLK(clk), .Q(\RF[15][10] ) );
  DFFPOSX1 \RF_reg[15][9]  ( .D(n3228), .CLK(clk), .Q(\RF[15][9] ) );
  DFFPOSX1 \RF_reg[15][8]  ( .D(n3227), .CLK(clk), .Q(\RF[15][8] ) );
  DFFPOSX1 \RF_reg[15][7]  ( .D(n3226), .CLK(clk), .Q(\RF[15][7] ) );
  DFFPOSX1 \RF_reg[15][6]  ( .D(n3225), .CLK(clk), .Q(\RF[15][6] ) );
  DFFPOSX1 \RF_reg[15][5]  ( .D(n3224), .CLK(clk), .Q(\RF[15][5] ) );
  DFFPOSX1 \RF_reg[15][4]  ( .D(n3223), .CLK(clk), .Q(\RF[15][4] ) );
  DFFPOSX1 \RF_reg[15][3]  ( .D(n3222), .CLK(clk), .Q(\RF[15][3] ) );
  DFFPOSX1 \RF_reg[15][2]  ( .D(n3221), .CLK(clk), .Q(\RF[15][2] ) );
  DFFPOSX1 \RF_reg[15][1]  ( .D(n3220), .CLK(clk), .Q(\RF[15][1] ) );
  DFFPOSX1 \RF_reg[15][0]  ( .D(n3219), .CLK(clk), .Q(\RF[15][0] ) );
  DFFPOSX1 \RF_reg[16][63]  ( .D(n3218), .CLK(clk), .Q(\RF[16][63] ) );
  DFFPOSX1 \RF_reg[16][62]  ( .D(n3217), .CLK(clk), .Q(\RF[16][62] ) );
  DFFPOSX1 \RF_reg[16][61]  ( .D(n3216), .CLK(clk), .Q(\RF[16][61] ) );
  DFFPOSX1 \RF_reg[16][60]  ( .D(n3215), .CLK(clk), .Q(\RF[16][60] ) );
  DFFPOSX1 \RF_reg[16][59]  ( .D(n3214), .CLK(clk), .Q(\RF[16][59] ) );
  DFFPOSX1 \RF_reg[16][58]  ( .D(n3213), .CLK(clk), .Q(\RF[16][58] ) );
  DFFPOSX1 \RF_reg[16][57]  ( .D(n3212), .CLK(clk), .Q(\RF[16][57] ) );
  DFFPOSX1 \RF_reg[16][56]  ( .D(n3211), .CLK(clk), .Q(\RF[16][56] ) );
  DFFPOSX1 \RF_reg[16][55]  ( .D(n3210), .CLK(clk), .Q(\RF[16][55] ) );
  DFFPOSX1 \RF_reg[16][54]  ( .D(n3209), .CLK(clk), .Q(\RF[16][54] ) );
  DFFPOSX1 \RF_reg[16][53]  ( .D(n3208), .CLK(clk), .Q(\RF[16][53] ) );
  DFFPOSX1 \RF_reg[16][52]  ( .D(n3207), .CLK(clk), .Q(\RF[16][52] ) );
  DFFPOSX1 \RF_reg[16][51]  ( .D(n3206), .CLK(clk), .Q(\RF[16][51] ) );
  DFFPOSX1 \RF_reg[16][50]  ( .D(n3205), .CLK(clk), .Q(\RF[16][50] ) );
  DFFPOSX1 \RF_reg[16][49]  ( .D(n3204), .CLK(clk), .Q(\RF[16][49] ) );
  DFFPOSX1 \RF_reg[16][48]  ( .D(n3203), .CLK(clk), .Q(\RF[16][48] ) );
  DFFPOSX1 \RF_reg[16][47]  ( .D(n3202), .CLK(clk), .Q(\RF[16][47] ) );
  DFFPOSX1 \RF_reg[16][46]  ( .D(n3201), .CLK(clk), .Q(\RF[16][46] ) );
  DFFPOSX1 \RF_reg[16][45]  ( .D(n3200), .CLK(clk), .Q(\RF[16][45] ) );
  DFFPOSX1 \RF_reg[16][44]  ( .D(n3199), .CLK(clk), .Q(\RF[16][44] ) );
  DFFPOSX1 \RF_reg[16][43]  ( .D(n3198), .CLK(clk), .Q(\RF[16][43] ) );
  DFFPOSX1 \RF_reg[16][42]  ( .D(n3197), .CLK(clk), .Q(\RF[16][42] ) );
  DFFPOSX1 \RF_reg[16][41]  ( .D(n3196), .CLK(clk), .Q(\RF[16][41] ) );
  DFFPOSX1 \RF_reg[16][40]  ( .D(n3195), .CLK(clk), .Q(\RF[16][40] ) );
  DFFPOSX1 \RF_reg[16][39]  ( .D(n3194), .CLK(clk), .Q(\RF[16][39] ) );
  DFFPOSX1 \RF_reg[16][38]  ( .D(n3193), .CLK(clk), .Q(\RF[16][38] ) );
  DFFPOSX1 \RF_reg[16][37]  ( .D(n3192), .CLK(clk), .Q(\RF[16][37] ) );
  DFFPOSX1 \RF_reg[16][36]  ( .D(n3191), .CLK(clk), .Q(\RF[16][36] ) );
  DFFPOSX1 \RF_reg[16][35]  ( .D(n3190), .CLK(clk), .Q(\RF[16][35] ) );
  DFFPOSX1 \RF_reg[16][34]  ( .D(n3189), .CLK(clk), .Q(\RF[16][34] ) );
  DFFPOSX1 \RF_reg[16][33]  ( .D(n3188), .CLK(clk), .Q(\RF[16][33] ) );
  DFFPOSX1 \RF_reg[16][32]  ( .D(n3187), .CLK(clk), .Q(\RF[16][32] ) );
  DFFPOSX1 \RF_reg[16][31]  ( .D(n3186), .CLK(clk), .Q(\RF[16][31] ) );
  DFFPOSX1 \RF_reg[16][30]  ( .D(n3185), .CLK(clk), .Q(\RF[16][30] ) );
  DFFPOSX1 \RF_reg[16][29]  ( .D(n3184), .CLK(clk), .Q(\RF[16][29] ) );
  DFFPOSX1 \RF_reg[16][28]  ( .D(n3183), .CLK(clk), .Q(\RF[16][28] ) );
  DFFPOSX1 \RF_reg[16][27]  ( .D(n3182), .CLK(clk), .Q(\RF[16][27] ) );
  DFFPOSX1 \RF_reg[16][26]  ( .D(n3181), .CLK(clk), .Q(\RF[16][26] ) );
  DFFPOSX1 \RF_reg[16][25]  ( .D(n3180), .CLK(clk), .Q(\RF[16][25] ) );
  DFFPOSX1 \RF_reg[16][24]  ( .D(n3179), .CLK(clk), .Q(\RF[16][24] ) );
  DFFPOSX1 \RF_reg[16][23]  ( .D(n3178), .CLK(clk), .Q(\RF[16][23] ) );
  DFFPOSX1 \RF_reg[16][22]  ( .D(n3177), .CLK(clk), .Q(\RF[16][22] ) );
  DFFPOSX1 \RF_reg[16][21]  ( .D(n3176), .CLK(clk), .Q(\RF[16][21] ) );
  DFFPOSX1 \RF_reg[16][20]  ( .D(n3175), .CLK(clk), .Q(\RF[16][20] ) );
  DFFPOSX1 \RF_reg[16][19]  ( .D(n3174), .CLK(clk), .Q(\RF[16][19] ) );
  DFFPOSX1 \RF_reg[16][18]  ( .D(n3173), .CLK(clk), .Q(\RF[16][18] ) );
  DFFPOSX1 \RF_reg[16][17]  ( .D(n3172), .CLK(clk), .Q(\RF[16][17] ) );
  DFFPOSX1 \RF_reg[16][16]  ( .D(n3171), .CLK(clk), .Q(\RF[16][16] ) );
  DFFPOSX1 \RF_reg[16][15]  ( .D(n3170), .CLK(clk), .Q(\RF[16][15] ) );
  DFFPOSX1 \RF_reg[16][14]  ( .D(n3169), .CLK(clk), .Q(\RF[16][14] ) );
  DFFPOSX1 \RF_reg[16][13]  ( .D(n3168), .CLK(clk), .Q(\RF[16][13] ) );
  DFFPOSX1 \RF_reg[16][12]  ( .D(n3167), .CLK(clk), .Q(\RF[16][12] ) );
  DFFPOSX1 \RF_reg[16][11]  ( .D(n3166), .CLK(clk), .Q(\RF[16][11] ) );
  DFFPOSX1 \RF_reg[16][10]  ( .D(n3165), .CLK(clk), .Q(\RF[16][10] ) );
  DFFPOSX1 \RF_reg[16][9]  ( .D(n3164), .CLK(clk), .Q(\RF[16][9] ) );
  DFFPOSX1 \RF_reg[16][8]  ( .D(n3163), .CLK(clk), .Q(\RF[16][8] ) );
  DFFPOSX1 \RF_reg[16][7]  ( .D(n3162), .CLK(clk), .Q(\RF[16][7] ) );
  DFFPOSX1 \RF_reg[16][6]  ( .D(n3161), .CLK(clk), .Q(\RF[16][6] ) );
  DFFPOSX1 \RF_reg[16][5]  ( .D(n3160), .CLK(clk), .Q(\RF[16][5] ) );
  DFFPOSX1 \RF_reg[16][4]  ( .D(n3159), .CLK(clk), .Q(\RF[16][4] ) );
  DFFPOSX1 \RF_reg[16][3]  ( .D(n3158), .CLK(clk), .Q(\RF[16][3] ) );
  DFFPOSX1 \RF_reg[16][2]  ( .D(n3157), .CLK(clk), .Q(\RF[16][2] ) );
  DFFPOSX1 \RF_reg[16][1]  ( .D(n3156), .CLK(clk), .Q(\RF[16][1] ) );
  DFFPOSX1 \RF_reg[16][0]  ( .D(n3155), .CLK(clk), .Q(\RF[16][0] ) );
  DFFPOSX1 \RF_reg[17][63]  ( .D(n3154), .CLK(clk), .Q(\RF[17][63] ) );
  DFFPOSX1 \RF_reg[17][62]  ( .D(n3153), .CLK(clk), .Q(\RF[17][62] ) );
  DFFPOSX1 \RF_reg[17][61]  ( .D(n3152), .CLK(clk), .Q(\RF[17][61] ) );
  DFFPOSX1 \RF_reg[17][60]  ( .D(n3151), .CLK(clk), .Q(\RF[17][60] ) );
  DFFPOSX1 \RF_reg[17][59]  ( .D(n3150), .CLK(clk), .Q(\RF[17][59] ) );
  DFFPOSX1 \RF_reg[17][58]  ( .D(n3149), .CLK(clk), .Q(\RF[17][58] ) );
  DFFPOSX1 \RF_reg[17][57]  ( .D(n3148), .CLK(clk), .Q(\RF[17][57] ) );
  DFFPOSX1 \RF_reg[17][56]  ( .D(n3147), .CLK(clk), .Q(\RF[17][56] ) );
  DFFPOSX1 \RF_reg[17][55]  ( .D(n3146), .CLK(clk), .Q(\RF[17][55] ) );
  DFFPOSX1 \RF_reg[17][54]  ( .D(n3145), .CLK(clk), .Q(\RF[17][54] ) );
  DFFPOSX1 \RF_reg[17][53]  ( .D(n3144), .CLK(clk), .Q(\RF[17][53] ) );
  DFFPOSX1 \RF_reg[17][52]  ( .D(n3143), .CLK(clk), .Q(\RF[17][52] ) );
  DFFPOSX1 \RF_reg[17][51]  ( .D(n3142), .CLK(clk), .Q(\RF[17][51] ) );
  DFFPOSX1 \RF_reg[17][50]  ( .D(n3141), .CLK(clk), .Q(\RF[17][50] ) );
  DFFPOSX1 \RF_reg[17][49]  ( .D(n3140), .CLK(clk), .Q(\RF[17][49] ) );
  DFFPOSX1 \RF_reg[17][48]  ( .D(n3139), .CLK(clk), .Q(\RF[17][48] ) );
  DFFPOSX1 \RF_reg[17][47]  ( .D(n3138), .CLK(clk), .Q(\RF[17][47] ) );
  DFFPOSX1 \RF_reg[17][46]  ( .D(n3137), .CLK(clk), .Q(\RF[17][46] ) );
  DFFPOSX1 \RF_reg[17][45]  ( .D(n3136), .CLK(clk), .Q(\RF[17][45] ) );
  DFFPOSX1 \RF_reg[17][44]  ( .D(n3135), .CLK(clk), .Q(\RF[17][44] ) );
  DFFPOSX1 \RF_reg[17][43]  ( .D(n3134), .CLK(clk), .Q(\RF[17][43] ) );
  DFFPOSX1 \RF_reg[17][42]  ( .D(n3133), .CLK(clk), .Q(\RF[17][42] ) );
  DFFPOSX1 \RF_reg[17][41]  ( .D(n3132), .CLK(clk), .Q(\RF[17][41] ) );
  DFFPOSX1 \RF_reg[17][40]  ( .D(n3131), .CLK(clk), .Q(\RF[17][40] ) );
  DFFPOSX1 \RF_reg[17][39]  ( .D(n3130), .CLK(clk), .Q(\RF[17][39] ) );
  DFFPOSX1 \RF_reg[17][38]  ( .D(n3129), .CLK(clk), .Q(\RF[17][38] ) );
  DFFPOSX1 \RF_reg[17][37]  ( .D(n3128), .CLK(clk), .Q(\RF[17][37] ) );
  DFFPOSX1 \RF_reg[17][36]  ( .D(n3127), .CLK(clk), .Q(\RF[17][36] ) );
  DFFPOSX1 \RF_reg[17][35]  ( .D(n3126), .CLK(clk), .Q(\RF[17][35] ) );
  DFFPOSX1 \RF_reg[17][34]  ( .D(n3125), .CLK(clk), .Q(\RF[17][34] ) );
  DFFPOSX1 \RF_reg[17][33]  ( .D(n3124), .CLK(clk), .Q(\RF[17][33] ) );
  DFFPOSX1 \RF_reg[17][32]  ( .D(n3123), .CLK(clk), .Q(\RF[17][32] ) );
  DFFPOSX1 \RF_reg[17][31]  ( .D(n3122), .CLK(clk), .Q(\RF[17][31] ) );
  DFFPOSX1 \RF_reg[17][30]  ( .D(n3121), .CLK(clk), .Q(\RF[17][30] ) );
  DFFPOSX1 \RF_reg[17][29]  ( .D(n3120), .CLK(clk), .Q(\RF[17][29] ) );
  DFFPOSX1 \RF_reg[17][28]  ( .D(n3119), .CLK(clk), .Q(\RF[17][28] ) );
  DFFPOSX1 \RF_reg[17][27]  ( .D(n3118), .CLK(clk), .Q(\RF[17][27] ) );
  DFFPOSX1 \RF_reg[17][26]  ( .D(n3117), .CLK(clk), .Q(\RF[17][26] ) );
  DFFPOSX1 \RF_reg[17][25]  ( .D(n3116), .CLK(clk), .Q(\RF[17][25] ) );
  DFFPOSX1 \RF_reg[17][24]  ( .D(n3115), .CLK(clk), .Q(\RF[17][24] ) );
  DFFPOSX1 \RF_reg[17][23]  ( .D(n3114), .CLK(clk), .Q(\RF[17][23] ) );
  DFFPOSX1 \RF_reg[17][22]  ( .D(n3113), .CLK(clk), .Q(\RF[17][22] ) );
  DFFPOSX1 \RF_reg[17][21]  ( .D(n3112), .CLK(clk), .Q(\RF[17][21] ) );
  DFFPOSX1 \RF_reg[17][20]  ( .D(n3111), .CLK(clk), .Q(\RF[17][20] ) );
  DFFPOSX1 \RF_reg[17][19]  ( .D(n3110), .CLK(clk), .Q(\RF[17][19] ) );
  DFFPOSX1 \RF_reg[17][18]  ( .D(n3109), .CLK(clk), .Q(\RF[17][18] ) );
  DFFPOSX1 \RF_reg[17][17]  ( .D(n3108), .CLK(clk), .Q(\RF[17][17] ) );
  DFFPOSX1 \RF_reg[17][16]  ( .D(n3107), .CLK(clk), .Q(\RF[17][16] ) );
  DFFPOSX1 \RF_reg[17][15]  ( .D(n3106), .CLK(clk), .Q(\RF[17][15] ) );
  DFFPOSX1 \RF_reg[17][14]  ( .D(n3105), .CLK(clk), .Q(\RF[17][14] ) );
  DFFPOSX1 \RF_reg[17][13]  ( .D(n3104), .CLK(clk), .Q(\RF[17][13] ) );
  DFFPOSX1 \RF_reg[17][12]  ( .D(n3103), .CLK(clk), .Q(\RF[17][12] ) );
  DFFPOSX1 \RF_reg[17][11]  ( .D(n3102), .CLK(clk), .Q(\RF[17][11] ) );
  DFFPOSX1 \RF_reg[17][10]  ( .D(n3101), .CLK(clk), .Q(\RF[17][10] ) );
  DFFPOSX1 \RF_reg[17][9]  ( .D(n3100), .CLK(clk), .Q(\RF[17][9] ) );
  DFFPOSX1 \RF_reg[17][8]  ( .D(n3099), .CLK(clk), .Q(\RF[17][8] ) );
  DFFPOSX1 \RF_reg[17][7]  ( .D(n3098), .CLK(clk), .Q(\RF[17][7] ) );
  DFFPOSX1 \RF_reg[17][6]  ( .D(n3097), .CLK(clk), .Q(\RF[17][6] ) );
  DFFPOSX1 \RF_reg[17][5]  ( .D(n3096), .CLK(clk), .Q(\RF[17][5] ) );
  DFFPOSX1 \RF_reg[17][4]  ( .D(n3095), .CLK(clk), .Q(\RF[17][4] ) );
  DFFPOSX1 \RF_reg[17][3]  ( .D(n3094), .CLK(clk), .Q(\RF[17][3] ) );
  DFFPOSX1 \RF_reg[17][2]  ( .D(n3093), .CLK(clk), .Q(\RF[17][2] ) );
  DFFPOSX1 \RF_reg[17][1]  ( .D(n3092), .CLK(clk), .Q(\RF[17][1] ) );
  DFFPOSX1 \RF_reg[17][0]  ( .D(n3091), .CLK(clk), .Q(\RF[17][0] ) );
  DFFPOSX1 \RF_reg[18][63]  ( .D(n3090), .CLK(clk), .Q(\RF[18][63] ) );
  DFFPOSX1 \RF_reg[18][62]  ( .D(n3089), .CLK(clk), .Q(\RF[18][62] ) );
  DFFPOSX1 \RF_reg[18][61]  ( .D(n3088), .CLK(clk), .Q(\RF[18][61] ) );
  DFFPOSX1 \RF_reg[18][60]  ( .D(n3087), .CLK(clk), .Q(\RF[18][60] ) );
  DFFPOSX1 \RF_reg[18][59]  ( .D(n3086), .CLK(clk), .Q(\RF[18][59] ) );
  DFFPOSX1 \RF_reg[18][58]  ( .D(n3085), .CLK(clk), .Q(\RF[18][58] ) );
  DFFPOSX1 \RF_reg[18][57]  ( .D(n3084), .CLK(clk), .Q(\RF[18][57] ) );
  DFFPOSX1 \RF_reg[18][56]  ( .D(n3083), .CLK(clk), .Q(\RF[18][56] ) );
  DFFPOSX1 \RF_reg[18][55]  ( .D(n3082), .CLK(clk), .Q(\RF[18][55] ) );
  DFFPOSX1 \RF_reg[18][54]  ( .D(n3081), .CLK(clk), .Q(\RF[18][54] ) );
  DFFPOSX1 \RF_reg[18][53]  ( .D(n3080), .CLK(clk), .Q(\RF[18][53] ) );
  DFFPOSX1 \RF_reg[18][52]  ( .D(n3079), .CLK(clk), .Q(\RF[18][52] ) );
  DFFPOSX1 \RF_reg[18][51]  ( .D(n3078), .CLK(clk), .Q(\RF[18][51] ) );
  DFFPOSX1 \RF_reg[18][50]  ( .D(n3077), .CLK(clk), .Q(\RF[18][50] ) );
  DFFPOSX1 \RF_reg[18][49]  ( .D(n3076), .CLK(clk), .Q(\RF[18][49] ) );
  DFFPOSX1 \RF_reg[18][48]  ( .D(n3075), .CLK(clk), .Q(\RF[18][48] ) );
  DFFPOSX1 \RF_reg[18][47]  ( .D(n3074), .CLK(clk), .Q(\RF[18][47] ) );
  DFFPOSX1 \RF_reg[18][46]  ( .D(n3073), .CLK(clk), .Q(\RF[18][46] ) );
  DFFPOSX1 \RF_reg[18][45]  ( .D(n3072), .CLK(clk), .Q(\RF[18][45] ) );
  DFFPOSX1 \RF_reg[18][44]  ( .D(n3071), .CLK(clk), .Q(\RF[18][44] ) );
  DFFPOSX1 \RF_reg[18][43]  ( .D(n3070), .CLK(clk), .Q(\RF[18][43] ) );
  DFFPOSX1 \RF_reg[18][42]  ( .D(n3069), .CLK(clk), .Q(\RF[18][42] ) );
  DFFPOSX1 \RF_reg[18][41]  ( .D(n3068), .CLK(clk), .Q(\RF[18][41] ) );
  DFFPOSX1 \RF_reg[18][40]  ( .D(n3067), .CLK(clk), .Q(\RF[18][40] ) );
  DFFPOSX1 \RF_reg[18][39]  ( .D(n3066), .CLK(clk), .Q(\RF[18][39] ) );
  DFFPOSX1 \RF_reg[18][38]  ( .D(n3065), .CLK(clk), .Q(\RF[18][38] ) );
  DFFPOSX1 \RF_reg[18][37]  ( .D(n3064), .CLK(clk), .Q(\RF[18][37] ) );
  DFFPOSX1 \RF_reg[18][36]  ( .D(n3063), .CLK(clk), .Q(\RF[18][36] ) );
  DFFPOSX1 \RF_reg[18][35]  ( .D(n3062), .CLK(clk), .Q(\RF[18][35] ) );
  DFFPOSX1 \RF_reg[18][34]  ( .D(n3061), .CLK(clk), .Q(\RF[18][34] ) );
  DFFPOSX1 \RF_reg[18][33]  ( .D(n3060), .CLK(clk), .Q(\RF[18][33] ) );
  DFFPOSX1 \RF_reg[18][32]  ( .D(n3059), .CLK(clk), .Q(\RF[18][32] ) );
  DFFPOSX1 \RF_reg[18][31]  ( .D(n3058), .CLK(clk), .Q(\RF[18][31] ) );
  DFFPOSX1 \RF_reg[18][30]  ( .D(n3057), .CLK(clk), .Q(\RF[18][30] ) );
  DFFPOSX1 \RF_reg[18][29]  ( .D(n3056), .CLK(clk), .Q(\RF[18][29] ) );
  DFFPOSX1 \RF_reg[18][28]  ( .D(n3055), .CLK(clk), .Q(\RF[18][28] ) );
  DFFPOSX1 \RF_reg[18][27]  ( .D(n3054), .CLK(clk), .Q(\RF[18][27] ) );
  DFFPOSX1 \RF_reg[18][26]  ( .D(n3053), .CLK(clk), .Q(\RF[18][26] ) );
  DFFPOSX1 \RF_reg[18][25]  ( .D(n3052), .CLK(clk), .Q(\RF[18][25] ) );
  DFFPOSX1 \RF_reg[18][24]  ( .D(n3051), .CLK(clk), .Q(\RF[18][24] ) );
  DFFPOSX1 \RF_reg[18][23]  ( .D(n3050), .CLK(clk), .Q(\RF[18][23] ) );
  DFFPOSX1 \RF_reg[18][22]  ( .D(n3049), .CLK(clk), .Q(\RF[18][22] ) );
  DFFPOSX1 \RF_reg[18][21]  ( .D(n3048), .CLK(clk), .Q(\RF[18][21] ) );
  DFFPOSX1 \RF_reg[18][20]  ( .D(n3047), .CLK(clk), .Q(\RF[18][20] ) );
  DFFPOSX1 \RF_reg[18][19]  ( .D(n3046), .CLK(clk), .Q(\RF[18][19] ) );
  DFFPOSX1 \RF_reg[18][18]  ( .D(n3045), .CLK(clk), .Q(\RF[18][18] ) );
  DFFPOSX1 \RF_reg[18][17]  ( .D(n3044), .CLK(clk), .Q(\RF[18][17] ) );
  DFFPOSX1 \RF_reg[18][16]  ( .D(n3043), .CLK(clk), .Q(\RF[18][16] ) );
  DFFPOSX1 \RF_reg[18][15]  ( .D(n3042), .CLK(clk), .Q(\RF[18][15] ) );
  DFFPOSX1 \RF_reg[18][14]  ( .D(n3041), .CLK(clk), .Q(\RF[18][14] ) );
  DFFPOSX1 \RF_reg[18][13]  ( .D(n3040), .CLK(clk), .Q(\RF[18][13] ) );
  DFFPOSX1 \RF_reg[18][12]  ( .D(n3039), .CLK(clk), .Q(\RF[18][12] ) );
  DFFPOSX1 \RF_reg[18][11]  ( .D(n3038), .CLK(clk), .Q(\RF[18][11] ) );
  DFFPOSX1 \RF_reg[18][10]  ( .D(n3037), .CLK(clk), .Q(\RF[18][10] ) );
  DFFPOSX1 \RF_reg[18][9]  ( .D(n3036), .CLK(clk), .Q(\RF[18][9] ) );
  DFFPOSX1 \RF_reg[18][8]  ( .D(n3035), .CLK(clk), .Q(\RF[18][8] ) );
  DFFPOSX1 \RF_reg[18][7]  ( .D(n3034), .CLK(clk), .Q(\RF[18][7] ) );
  DFFPOSX1 \RF_reg[18][6]  ( .D(n3033), .CLK(clk), .Q(\RF[18][6] ) );
  DFFPOSX1 \RF_reg[18][5]  ( .D(n3032), .CLK(clk), .Q(\RF[18][5] ) );
  DFFPOSX1 \RF_reg[18][4]  ( .D(n3031), .CLK(clk), .Q(\RF[18][4] ) );
  DFFPOSX1 \RF_reg[18][3]  ( .D(n3030), .CLK(clk), .Q(\RF[18][3] ) );
  DFFPOSX1 \RF_reg[18][2]  ( .D(n3029), .CLK(clk), .Q(\RF[18][2] ) );
  DFFPOSX1 \RF_reg[18][1]  ( .D(n3028), .CLK(clk), .Q(\RF[18][1] ) );
  DFFPOSX1 \RF_reg[18][0]  ( .D(n3027), .CLK(clk), .Q(\RF[18][0] ) );
  DFFPOSX1 \RF_reg[19][63]  ( .D(n3026), .CLK(clk), .Q(\RF[19][63] ) );
  DFFPOSX1 \RF_reg[19][62]  ( .D(n3025), .CLK(clk), .Q(\RF[19][62] ) );
  DFFPOSX1 \RF_reg[19][61]  ( .D(n3024), .CLK(clk), .Q(\RF[19][61] ) );
  DFFPOSX1 \RF_reg[19][60]  ( .D(n3023), .CLK(clk), .Q(\RF[19][60] ) );
  DFFPOSX1 \RF_reg[19][59]  ( .D(n3022), .CLK(clk), .Q(\RF[19][59] ) );
  DFFPOSX1 \RF_reg[19][58]  ( .D(n3021), .CLK(clk), .Q(\RF[19][58] ) );
  DFFPOSX1 \RF_reg[19][57]  ( .D(n3020), .CLK(clk), .Q(\RF[19][57] ) );
  DFFPOSX1 \RF_reg[19][56]  ( .D(n3019), .CLK(clk), .Q(\RF[19][56] ) );
  DFFPOSX1 \RF_reg[19][55]  ( .D(n3018), .CLK(clk), .Q(\RF[19][55] ) );
  DFFPOSX1 \RF_reg[19][54]  ( .D(n3017), .CLK(clk), .Q(\RF[19][54] ) );
  DFFPOSX1 \RF_reg[19][53]  ( .D(n3016), .CLK(clk), .Q(\RF[19][53] ) );
  DFFPOSX1 \RF_reg[19][52]  ( .D(n3015), .CLK(clk), .Q(\RF[19][52] ) );
  DFFPOSX1 \RF_reg[19][51]  ( .D(n3014), .CLK(clk), .Q(\RF[19][51] ) );
  DFFPOSX1 \RF_reg[19][50]  ( .D(n3013), .CLK(clk), .Q(\RF[19][50] ) );
  DFFPOSX1 \RF_reg[19][49]  ( .D(n3012), .CLK(clk), .Q(\RF[19][49] ) );
  DFFPOSX1 \RF_reg[19][48]  ( .D(n3011), .CLK(clk), .Q(\RF[19][48] ) );
  DFFPOSX1 \RF_reg[19][47]  ( .D(n3010), .CLK(clk), .Q(\RF[19][47] ) );
  DFFPOSX1 \RF_reg[19][46]  ( .D(n3009), .CLK(clk), .Q(\RF[19][46] ) );
  DFFPOSX1 \RF_reg[19][45]  ( .D(n3008), .CLK(clk), .Q(\RF[19][45] ) );
  DFFPOSX1 \RF_reg[19][44]  ( .D(n3007), .CLK(clk), .Q(\RF[19][44] ) );
  DFFPOSX1 \RF_reg[19][43]  ( .D(n3006), .CLK(clk), .Q(\RF[19][43] ) );
  DFFPOSX1 \RF_reg[19][42]  ( .D(n3005), .CLK(clk), .Q(\RF[19][42] ) );
  DFFPOSX1 \RF_reg[19][41]  ( .D(n3004), .CLK(clk), .Q(\RF[19][41] ) );
  DFFPOSX1 \RF_reg[19][40]  ( .D(n3003), .CLK(clk), .Q(\RF[19][40] ) );
  DFFPOSX1 \RF_reg[19][39]  ( .D(n3002), .CLK(clk), .Q(\RF[19][39] ) );
  DFFPOSX1 \RF_reg[19][38]  ( .D(n3001), .CLK(clk), .Q(\RF[19][38] ) );
  DFFPOSX1 \RF_reg[19][37]  ( .D(n3000), .CLK(clk), .Q(\RF[19][37] ) );
  DFFPOSX1 \RF_reg[19][36]  ( .D(n2999), .CLK(clk), .Q(\RF[19][36] ) );
  DFFPOSX1 \RF_reg[19][35]  ( .D(n2998), .CLK(clk), .Q(\RF[19][35] ) );
  DFFPOSX1 \RF_reg[19][34]  ( .D(n2997), .CLK(clk), .Q(\RF[19][34] ) );
  DFFPOSX1 \RF_reg[19][33]  ( .D(n2996), .CLK(clk), .Q(\RF[19][33] ) );
  DFFPOSX1 \RF_reg[19][32]  ( .D(n2995), .CLK(clk), .Q(\RF[19][32] ) );
  DFFPOSX1 \RF_reg[19][31]  ( .D(n2994), .CLK(clk), .Q(\RF[19][31] ) );
  DFFPOSX1 \RF_reg[19][30]  ( .D(n2993), .CLK(clk), .Q(\RF[19][30] ) );
  DFFPOSX1 \RF_reg[19][29]  ( .D(n2992), .CLK(clk), .Q(\RF[19][29] ) );
  DFFPOSX1 \RF_reg[19][28]  ( .D(n2991), .CLK(clk), .Q(\RF[19][28] ) );
  DFFPOSX1 \RF_reg[19][27]  ( .D(n2990), .CLK(clk), .Q(\RF[19][27] ) );
  DFFPOSX1 \RF_reg[19][26]  ( .D(n2989), .CLK(clk), .Q(\RF[19][26] ) );
  DFFPOSX1 \RF_reg[19][25]  ( .D(n2988), .CLK(clk), .Q(\RF[19][25] ) );
  DFFPOSX1 \RF_reg[19][24]  ( .D(n2987), .CLK(clk), .Q(\RF[19][24] ) );
  DFFPOSX1 \RF_reg[19][23]  ( .D(n2986), .CLK(clk), .Q(\RF[19][23] ) );
  DFFPOSX1 \RF_reg[19][22]  ( .D(n2985), .CLK(clk), .Q(\RF[19][22] ) );
  DFFPOSX1 \RF_reg[19][21]  ( .D(n2984), .CLK(clk), .Q(\RF[19][21] ) );
  DFFPOSX1 \RF_reg[19][20]  ( .D(n2983), .CLK(clk), .Q(\RF[19][20] ) );
  DFFPOSX1 \RF_reg[19][19]  ( .D(n2982), .CLK(clk), .Q(\RF[19][19] ) );
  DFFPOSX1 \RF_reg[19][18]  ( .D(n2981), .CLK(clk), .Q(\RF[19][18] ) );
  DFFPOSX1 \RF_reg[19][17]  ( .D(n2980), .CLK(clk), .Q(\RF[19][17] ) );
  DFFPOSX1 \RF_reg[19][16]  ( .D(n2979), .CLK(clk), .Q(\RF[19][16] ) );
  DFFPOSX1 \RF_reg[19][15]  ( .D(n2978), .CLK(clk), .Q(\RF[19][15] ) );
  DFFPOSX1 \RF_reg[19][14]  ( .D(n2977), .CLK(clk), .Q(\RF[19][14] ) );
  DFFPOSX1 \RF_reg[19][13]  ( .D(n2976), .CLK(clk), .Q(\RF[19][13] ) );
  DFFPOSX1 \RF_reg[19][12]  ( .D(n2975), .CLK(clk), .Q(\RF[19][12] ) );
  DFFPOSX1 \RF_reg[19][11]  ( .D(n2974), .CLK(clk), .Q(\RF[19][11] ) );
  DFFPOSX1 \RF_reg[19][10]  ( .D(n2973), .CLK(clk), .Q(\RF[19][10] ) );
  DFFPOSX1 \RF_reg[19][9]  ( .D(n2972), .CLK(clk), .Q(\RF[19][9] ) );
  DFFPOSX1 \RF_reg[19][8]  ( .D(n2971), .CLK(clk), .Q(\RF[19][8] ) );
  DFFPOSX1 \RF_reg[19][7]  ( .D(n2970), .CLK(clk), .Q(\RF[19][7] ) );
  DFFPOSX1 \RF_reg[19][6]  ( .D(n2969), .CLK(clk), .Q(\RF[19][6] ) );
  DFFPOSX1 \RF_reg[19][5]  ( .D(n2968), .CLK(clk), .Q(\RF[19][5] ) );
  DFFPOSX1 \RF_reg[19][4]  ( .D(n2967), .CLK(clk), .Q(\RF[19][4] ) );
  DFFPOSX1 \RF_reg[19][3]  ( .D(n2966), .CLK(clk), .Q(\RF[19][3] ) );
  DFFPOSX1 \RF_reg[19][2]  ( .D(n2965), .CLK(clk), .Q(\RF[19][2] ) );
  DFFPOSX1 \RF_reg[19][1]  ( .D(n2964), .CLK(clk), .Q(\RF[19][1] ) );
  DFFPOSX1 \RF_reg[19][0]  ( .D(n2963), .CLK(clk), .Q(\RF[19][0] ) );
  DFFPOSX1 \RF_reg[20][63]  ( .D(n2962), .CLK(clk), .Q(\RF[20][63] ) );
  DFFPOSX1 \RF_reg[20][62]  ( .D(n2961), .CLK(clk), .Q(\RF[20][62] ) );
  DFFPOSX1 \RF_reg[20][61]  ( .D(n2960), .CLK(clk), .Q(\RF[20][61] ) );
  DFFPOSX1 \RF_reg[20][60]  ( .D(n2959), .CLK(clk), .Q(\RF[20][60] ) );
  DFFPOSX1 \RF_reg[20][59]  ( .D(n2958), .CLK(clk), .Q(\RF[20][59] ) );
  DFFPOSX1 \RF_reg[20][58]  ( .D(n2957), .CLK(clk), .Q(\RF[20][58] ) );
  DFFPOSX1 \RF_reg[20][57]  ( .D(n2956), .CLK(clk), .Q(\RF[20][57] ) );
  DFFPOSX1 \RF_reg[20][56]  ( .D(n2955), .CLK(clk), .Q(\RF[20][56] ) );
  DFFPOSX1 \RF_reg[20][55]  ( .D(n2954), .CLK(clk), .Q(\RF[20][55] ) );
  DFFPOSX1 \RF_reg[20][54]  ( .D(n2953), .CLK(clk), .Q(\RF[20][54] ) );
  DFFPOSX1 \RF_reg[20][53]  ( .D(n2952), .CLK(clk), .Q(\RF[20][53] ) );
  DFFPOSX1 \RF_reg[20][52]  ( .D(n2951), .CLK(clk), .Q(\RF[20][52] ) );
  DFFPOSX1 \RF_reg[20][51]  ( .D(n2950), .CLK(clk), .Q(\RF[20][51] ) );
  DFFPOSX1 \RF_reg[20][50]  ( .D(n2949), .CLK(clk), .Q(\RF[20][50] ) );
  DFFPOSX1 \RF_reg[20][49]  ( .D(n2948), .CLK(clk), .Q(\RF[20][49] ) );
  DFFPOSX1 \RF_reg[20][48]  ( .D(n2947), .CLK(clk), .Q(\RF[20][48] ) );
  DFFPOSX1 \RF_reg[20][47]  ( .D(n2946), .CLK(clk), .Q(\RF[20][47] ) );
  DFFPOSX1 \RF_reg[20][46]  ( .D(n2945), .CLK(clk), .Q(\RF[20][46] ) );
  DFFPOSX1 \RF_reg[20][45]  ( .D(n2944), .CLK(clk), .Q(\RF[20][45] ) );
  DFFPOSX1 \RF_reg[20][44]  ( .D(n2943), .CLK(clk), .Q(\RF[20][44] ) );
  DFFPOSX1 \RF_reg[20][43]  ( .D(n2942), .CLK(clk), .Q(\RF[20][43] ) );
  DFFPOSX1 \RF_reg[20][42]  ( .D(n2941), .CLK(clk), .Q(\RF[20][42] ) );
  DFFPOSX1 \RF_reg[20][41]  ( .D(n2940), .CLK(clk), .Q(\RF[20][41] ) );
  DFFPOSX1 \RF_reg[20][40]  ( .D(n2939), .CLK(clk), .Q(\RF[20][40] ) );
  DFFPOSX1 \RF_reg[20][39]  ( .D(n2938), .CLK(clk), .Q(\RF[20][39] ) );
  DFFPOSX1 \RF_reg[20][38]  ( .D(n2937), .CLK(clk), .Q(\RF[20][38] ) );
  DFFPOSX1 \RF_reg[20][37]  ( .D(n2936), .CLK(clk), .Q(\RF[20][37] ) );
  DFFPOSX1 \RF_reg[20][36]  ( .D(n2935), .CLK(clk), .Q(\RF[20][36] ) );
  DFFPOSX1 \RF_reg[20][35]  ( .D(n2934), .CLK(clk), .Q(\RF[20][35] ) );
  DFFPOSX1 \RF_reg[20][34]  ( .D(n2933), .CLK(clk), .Q(\RF[20][34] ) );
  DFFPOSX1 \RF_reg[20][33]  ( .D(n2932), .CLK(clk), .Q(\RF[20][33] ) );
  DFFPOSX1 \RF_reg[20][32]  ( .D(n2931), .CLK(clk), .Q(\RF[20][32] ) );
  DFFPOSX1 \RF_reg[20][31]  ( .D(n2930), .CLK(clk), .Q(\RF[20][31] ) );
  DFFPOSX1 \RF_reg[20][30]  ( .D(n2929), .CLK(clk), .Q(\RF[20][30] ) );
  DFFPOSX1 \RF_reg[20][29]  ( .D(n2928), .CLK(clk), .Q(\RF[20][29] ) );
  DFFPOSX1 \RF_reg[20][28]  ( .D(n2927), .CLK(clk), .Q(\RF[20][28] ) );
  DFFPOSX1 \RF_reg[20][27]  ( .D(n2926), .CLK(clk), .Q(\RF[20][27] ) );
  DFFPOSX1 \RF_reg[20][26]  ( .D(n2925), .CLK(clk), .Q(\RF[20][26] ) );
  DFFPOSX1 \RF_reg[20][25]  ( .D(n2924), .CLK(clk), .Q(\RF[20][25] ) );
  DFFPOSX1 \RF_reg[20][24]  ( .D(n2923), .CLK(clk), .Q(\RF[20][24] ) );
  DFFPOSX1 \RF_reg[20][23]  ( .D(n2922), .CLK(clk), .Q(\RF[20][23] ) );
  DFFPOSX1 \RF_reg[20][22]  ( .D(n2921), .CLK(clk), .Q(\RF[20][22] ) );
  DFFPOSX1 \RF_reg[20][21]  ( .D(n2920), .CLK(clk), .Q(\RF[20][21] ) );
  DFFPOSX1 \RF_reg[20][20]  ( .D(n2919), .CLK(clk), .Q(\RF[20][20] ) );
  DFFPOSX1 \RF_reg[20][19]  ( .D(n2918), .CLK(clk), .Q(\RF[20][19] ) );
  DFFPOSX1 \RF_reg[20][18]  ( .D(n2917), .CLK(clk), .Q(\RF[20][18] ) );
  DFFPOSX1 \RF_reg[20][17]  ( .D(n2916), .CLK(clk), .Q(\RF[20][17] ) );
  DFFPOSX1 \RF_reg[20][16]  ( .D(n2915), .CLK(clk), .Q(\RF[20][16] ) );
  DFFPOSX1 \RF_reg[20][15]  ( .D(n2914), .CLK(clk), .Q(\RF[20][15] ) );
  DFFPOSX1 \RF_reg[20][14]  ( .D(n2913), .CLK(clk), .Q(\RF[20][14] ) );
  DFFPOSX1 \RF_reg[20][13]  ( .D(n2912), .CLK(clk), .Q(\RF[20][13] ) );
  DFFPOSX1 \RF_reg[20][12]  ( .D(n2911), .CLK(clk), .Q(\RF[20][12] ) );
  DFFPOSX1 \RF_reg[20][11]  ( .D(n2910), .CLK(clk), .Q(\RF[20][11] ) );
  DFFPOSX1 \RF_reg[20][10]  ( .D(n2909), .CLK(clk), .Q(\RF[20][10] ) );
  DFFPOSX1 \RF_reg[20][9]  ( .D(n2908), .CLK(clk), .Q(\RF[20][9] ) );
  DFFPOSX1 \RF_reg[20][8]  ( .D(n2907), .CLK(clk), .Q(\RF[20][8] ) );
  DFFPOSX1 \RF_reg[20][7]  ( .D(n2906), .CLK(clk), .Q(\RF[20][7] ) );
  DFFPOSX1 \RF_reg[20][6]  ( .D(n2905), .CLK(clk), .Q(\RF[20][6] ) );
  DFFPOSX1 \RF_reg[20][5]  ( .D(n2904), .CLK(clk), .Q(\RF[20][5] ) );
  DFFPOSX1 \RF_reg[20][4]  ( .D(n2903), .CLK(clk), .Q(\RF[20][4] ) );
  DFFPOSX1 \RF_reg[20][3]  ( .D(n2902), .CLK(clk), .Q(\RF[20][3] ) );
  DFFPOSX1 \RF_reg[20][2]  ( .D(n2901), .CLK(clk), .Q(\RF[20][2] ) );
  DFFPOSX1 \RF_reg[20][1]  ( .D(n2900), .CLK(clk), .Q(\RF[20][1] ) );
  DFFPOSX1 \RF_reg[20][0]  ( .D(n2899), .CLK(clk), .Q(\RF[20][0] ) );
  DFFPOSX1 \RF_reg[21][63]  ( .D(n2898), .CLK(clk), .Q(\RF[21][63] ) );
  DFFPOSX1 \RF_reg[21][62]  ( .D(n2897), .CLK(clk), .Q(\RF[21][62] ) );
  DFFPOSX1 \RF_reg[21][61]  ( .D(n2896), .CLK(clk), .Q(\RF[21][61] ) );
  DFFPOSX1 \RF_reg[21][60]  ( .D(n2895), .CLK(clk), .Q(\RF[21][60] ) );
  DFFPOSX1 \RF_reg[21][59]  ( .D(n2894), .CLK(clk), .Q(\RF[21][59] ) );
  DFFPOSX1 \RF_reg[21][58]  ( .D(n2893), .CLK(clk), .Q(\RF[21][58] ) );
  DFFPOSX1 \RF_reg[21][57]  ( .D(n2892), .CLK(clk), .Q(\RF[21][57] ) );
  DFFPOSX1 \RF_reg[21][56]  ( .D(n2891), .CLK(clk), .Q(\RF[21][56] ) );
  DFFPOSX1 \RF_reg[21][55]  ( .D(n2890), .CLK(clk), .Q(\RF[21][55] ) );
  DFFPOSX1 \RF_reg[21][54]  ( .D(n2889), .CLK(clk), .Q(\RF[21][54] ) );
  DFFPOSX1 \RF_reg[21][53]  ( .D(n2888), .CLK(clk), .Q(\RF[21][53] ) );
  DFFPOSX1 \RF_reg[21][52]  ( .D(n2887), .CLK(clk), .Q(\RF[21][52] ) );
  DFFPOSX1 \RF_reg[21][51]  ( .D(n2886), .CLK(clk), .Q(\RF[21][51] ) );
  DFFPOSX1 \RF_reg[21][50]  ( .D(n2885), .CLK(clk), .Q(\RF[21][50] ) );
  DFFPOSX1 \RF_reg[21][49]  ( .D(n2884), .CLK(clk), .Q(\RF[21][49] ) );
  DFFPOSX1 \RF_reg[21][48]  ( .D(n2883), .CLK(clk), .Q(\RF[21][48] ) );
  DFFPOSX1 \RF_reg[21][47]  ( .D(n2882), .CLK(clk), .Q(\RF[21][47] ) );
  DFFPOSX1 \RF_reg[21][46]  ( .D(n2881), .CLK(clk), .Q(\RF[21][46] ) );
  DFFPOSX1 \RF_reg[21][45]  ( .D(n2880), .CLK(clk), .Q(\RF[21][45] ) );
  DFFPOSX1 \RF_reg[21][44]  ( .D(n2879), .CLK(clk), .Q(\RF[21][44] ) );
  DFFPOSX1 \RF_reg[21][43]  ( .D(n2878), .CLK(clk), .Q(\RF[21][43] ) );
  DFFPOSX1 \RF_reg[21][42]  ( .D(n2877), .CLK(clk), .Q(\RF[21][42] ) );
  DFFPOSX1 \RF_reg[21][41]  ( .D(n2876), .CLK(clk), .Q(\RF[21][41] ) );
  DFFPOSX1 \RF_reg[21][40]  ( .D(n2875), .CLK(clk), .Q(\RF[21][40] ) );
  DFFPOSX1 \RF_reg[21][39]  ( .D(n2874), .CLK(clk), .Q(\RF[21][39] ) );
  DFFPOSX1 \RF_reg[21][38]  ( .D(n2873), .CLK(clk), .Q(\RF[21][38] ) );
  DFFPOSX1 \RF_reg[21][37]  ( .D(n2872), .CLK(clk), .Q(\RF[21][37] ) );
  DFFPOSX1 \RF_reg[21][36]  ( .D(n2871), .CLK(clk), .Q(\RF[21][36] ) );
  DFFPOSX1 \RF_reg[21][35]  ( .D(n2870), .CLK(clk), .Q(\RF[21][35] ) );
  DFFPOSX1 \RF_reg[21][34]  ( .D(n2869), .CLK(clk), .Q(\RF[21][34] ) );
  DFFPOSX1 \RF_reg[21][33]  ( .D(n2868), .CLK(clk), .Q(\RF[21][33] ) );
  DFFPOSX1 \RF_reg[21][32]  ( .D(n2867), .CLK(clk), .Q(\RF[21][32] ) );
  DFFPOSX1 \RF_reg[21][31]  ( .D(n2866), .CLK(clk), .Q(\RF[21][31] ) );
  DFFPOSX1 \RF_reg[21][30]  ( .D(n2865), .CLK(clk), .Q(\RF[21][30] ) );
  DFFPOSX1 \RF_reg[21][29]  ( .D(n2864), .CLK(clk), .Q(\RF[21][29] ) );
  DFFPOSX1 \RF_reg[21][28]  ( .D(n2863), .CLK(clk), .Q(\RF[21][28] ) );
  DFFPOSX1 \RF_reg[21][27]  ( .D(n2862), .CLK(clk), .Q(\RF[21][27] ) );
  DFFPOSX1 \RF_reg[21][26]  ( .D(n2861), .CLK(clk), .Q(\RF[21][26] ) );
  DFFPOSX1 \RF_reg[21][25]  ( .D(n2860), .CLK(clk), .Q(\RF[21][25] ) );
  DFFPOSX1 \RF_reg[21][24]  ( .D(n2859), .CLK(clk), .Q(\RF[21][24] ) );
  DFFPOSX1 \RF_reg[21][23]  ( .D(n2858), .CLK(clk), .Q(\RF[21][23] ) );
  DFFPOSX1 \RF_reg[21][22]  ( .D(n2857), .CLK(clk), .Q(\RF[21][22] ) );
  DFFPOSX1 \RF_reg[21][21]  ( .D(n2856), .CLK(clk), .Q(\RF[21][21] ) );
  DFFPOSX1 \RF_reg[21][20]  ( .D(n2855), .CLK(clk), .Q(\RF[21][20] ) );
  DFFPOSX1 \RF_reg[21][19]  ( .D(n2854), .CLK(clk), .Q(\RF[21][19] ) );
  DFFPOSX1 \RF_reg[21][18]  ( .D(n2853), .CLK(clk), .Q(\RF[21][18] ) );
  DFFPOSX1 \RF_reg[21][17]  ( .D(n2852), .CLK(clk), .Q(\RF[21][17] ) );
  DFFPOSX1 \RF_reg[21][16]  ( .D(n2851), .CLK(clk), .Q(\RF[21][16] ) );
  DFFPOSX1 \RF_reg[21][15]  ( .D(n2850), .CLK(clk), .Q(\RF[21][15] ) );
  DFFPOSX1 \RF_reg[21][14]  ( .D(n2849), .CLK(clk), .Q(\RF[21][14] ) );
  DFFPOSX1 \RF_reg[21][13]  ( .D(n2848), .CLK(clk), .Q(\RF[21][13] ) );
  DFFPOSX1 \RF_reg[21][12]  ( .D(n2847), .CLK(clk), .Q(\RF[21][12] ) );
  DFFPOSX1 \RF_reg[21][11]  ( .D(n2846), .CLK(clk), .Q(\RF[21][11] ) );
  DFFPOSX1 \RF_reg[21][10]  ( .D(n2845), .CLK(clk), .Q(\RF[21][10] ) );
  DFFPOSX1 \RF_reg[21][9]  ( .D(n2844), .CLK(clk), .Q(\RF[21][9] ) );
  DFFPOSX1 \RF_reg[21][8]  ( .D(n2843), .CLK(clk), .Q(\RF[21][8] ) );
  DFFPOSX1 \RF_reg[21][7]  ( .D(n2842), .CLK(clk), .Q(\RF[21][7] ) );
  DFFPOSX1 \RF_reg[21][6]  ( .D(n2841), .CLK(clk), .Q(\RF[21][6] ) );
  DFFPOSX1 \RF_reg[21][5]  ( .D(n2840), .CLK(clk), .Q(\RF[21][5] ) );
  DFFPOSX1 \RF_reg[21][4]  ( .D(n2839), .CLK(clk), .Q(\RF[21][4] ) );
  DFFPOSX1 \RF_reg[21][3]  ( .D(n2838), .CLK(clk), .Q(\RF[21][3] ) );
  DFFPOSX1 \RF_reg[21][2]  ( .D(n2837), .CLK(clk), .Q(\RF[21][2] ) );
  DFFPOSX1 \RF_reg[21][1]  ( .D(n2836), .CLK(clk), .Q(\RF[21][1] ) );
  DFFPOSX1 \RF_reg[21][0]  ( .D(n2835), .CLK(clk), .Q(\RF[21][0] ) );
  DFFPOSX1 \RF_reg[22][63]  ( .D(n2834), .CLK(clk), .Q(\RF[22][63] ) );
  DFFPOSX1 \RF_reg[22][62]  ( .D(n2833), .CLK(clk), .Q(\RF[22][62] ) );
  DFFPOSX1 \RF_reg[22][61]  ( .D(n2832), .CLK(clk), .Q(\RF[22][61] ) );
  DFFPOSX1 \RF_reg[22][60]  ( .D(n2831), .CLK(clk), .Q(\RF[22][60] ) );
  DFFPOSX1 \RF_reg[22][59]  ( .D(n2830), .CLK(clk), .Q(\RF[22][59] ) );
  DFFPOSX1 \RF_reg[22][58]  ( .D(n2829), .CLK(clk), .Q(\RF[22][58] ) );
  DFFPOSX1 \RF_reg[22][57]  ( .D(n2828), .CLK(clk), .Q(\RF[22][57] ) );
  DFFPOSX1 \RF_reg[22][56]  ( .D(n2827), .CLK(clk), .Q(\RF[22][56] ) );
  DFFPOSX1 \RF_reg[22][55]  ( .D(n2826), .CLK(clk), .Q(\RF[22][55] ) );
  DFFPOSX1 \RF_reg[22][54]  ( .D(n2825), .CLK(clk), .Q(\RF[22][54] ) );
  DFFPOSX1 \RF_reg[22][53]  ( .D(n2824), .CLK(clk), .Q(\RF[22][53] ) );
  DFFPOSX1 \RF_reg[22][52]  ( .D(n2823), .CLK(clk), .Q(\RF[22][52] ) );
  DFFPOSX1 \RF_reg[22][51]  ( .D(n2822), .CLK(clk), .Q(\RF[22][51] ) );
  DFFPOSX1 \RF_reg[22][50]  ( .D(n2821), .CLK(clk), .Q(\RF[22][50] ) );
  DFFPOSX1 \RF_reg[22][49]  ( .D(n2820), .CLK(clk), .Q(\RF[22][49] ) );
  DFFPOSX1 \RF_reg[22][48]  ( .D(n2819), .CLK(clk), .Q(\RF[22][48] ) );
  DFFPOSX1 \RF_reg[22][47]  ( .D(n2818), .CLK(clk), .Q(\RF[22][47] ) );
  DFFPOSX1 \RF_reg[22][46]  ( .D(n2817), .CLK(clk), .Q(\RF[22][46] ) );
  DFFPOSX1 \RF_reg[22][45]  ( .D(n2816), .CLK(clk), .Q(\RF[22][45] ) );
  DFFPOSX1 \RF_reg[22][44]  ( .D(n2815), .CLK(clk), .Q(\RF[22][44] ) );
  DFFPOSX1 \RF_reg[22][43]  ( .D(n2814), .CLK(clk), .Q(\RF[22][43] ) );
  DFFPOSX1 \RF_reg[22][42]  ( .D(n2813), .CLK(clk), .Q(\RF[22][42] ) );
  DFFPOSX1 \RF_reg[22][41]  ( .D(n2812), .CLK(clk), .Q(\RF[22][41] ) );
  DFFPOSX1 \RF_reg[22][40]  ( .D(n2811), .CLK(clk), .Q(\RF[22][40] ) );
  DFFPOSX1 \RF_reg[22][39]  ( .D(n2810), .CLK(clk), .Q(\RF[22][39] ) );
  DFFPOSX1 \RF_reg[22][38]  ( .D(n2809), .CLK(clk), .Q(\RF[22][38] ) );
  DFFPOSX1 \RF_reg[22][37]  ( .D(n2808), .CLK(clk), .Q(\RF[22][37] ) );
  DFFPOSX1 \RF_reg[22][36]  ( .D(n2807), .CLK(clk), .Q(\RF[22][36] ) );
  DFFPOSX1 \RF_reg[22][35]  ( .D(n2806), .CLK(clk), .Q(\RF[22][35] ) );
  DFFPOSX1 \RF_reg[22][34]  ( .D(n2805), .CLK(clk), .Q(\RF[22][34] ) );
  DFFPOSX1 \RF_reg[22][33]  ( .D(n2804), .CLK(clk), .Q(\RF[22][33] ) );
  DFFPOSX1 \RF_reg[22][32]  ( .D(n2803), .CLK(clk), .Q(\RF[22][32] ) );
  DFFPOSX1 \RF_reg[22][31]  ( .D(n2802), .CLK(clk), .Q(\RF[22][31] ) );
  DFFPOSX1 \RF_reg[22][30]  ( .D(n2801), .CLK(clk), .Q(\RF[22][30] ) );
  DFFPOSX1 \RF_reg[22][29]  ( .D(n2800), .CLK(clk), .Q(\RF[22][29] ) );
  DFFPOSX1 \RF_reg[22][28]  ( .D(n2799), .CLK(clk), .Q(\RF[22][28] ) );
  DFFPOSX1 \RF_reg[22][27]  ( .D(n2798), .CLK(clk), .Q(\RF[22][27] ) );
  DFFPOSX1 \RF_reg[22][26]  ( .D(n2797), .CLK(clk), .Q(\RF[22][26] ) );
  DFFPOSX1 \RF_reg[22][25]  ( .D(n2796), .CLK(clk), .Q(\RF[22][25] ) );
  DFFPOSX1 \RF_reg[22][24]  ( .D(n2795), .CLK(clk), .Q(\RF[22][24] ) );
  DFFPOSX1 \RF_reg[22][23]  ( .D(n2794), .CLK(clk), .Q(\RF[22][23] ) );
  DFFPOSX1 \RF_reg[22][22]  ( .D(n2793), .CLK(clk), .Q(\RF[22][22] ) );
  DFFPOSX1 \RF_reg[22][21]  ( .D(n2792), .CLK(clk), .Q(\RF[22][21] ) );
  DFFPOSX1 \RF_reg[22][20]  ( .D(n2791), .CLK(clk), .Q(\RF[22][20] ) );
  DFFPOSX1 \RF_reg[22][19]  ( .D(n2790), .CLK(clk), .Q(\RF[22][19] ) );
  DFFPOSX1 \RF_reg[22][18]  ( .D(n2789), .CLK(clk), .Q(\RF[22][18] ) );
  DFFPOSX1 \RF_reg[22][17]  ( .D(n2788), .CLK(clk), .Q(\RF[22][17] ) );
  DFFPOSX1 \RF_reg[22][16]  ( .D(n2787), .CLK(clk), .Q(\RF[22][16] ) );
  DFFPOSX1 \RF_reg[22][15]  ( .D(n2786), .CLK(clk), .Q(\RF[22][15] ) );
  DFFPOSX1 \RF_reg[22][14]  ( .D(n2785), .CLK(clk), .Q(\RF[22][14] ) );
  DFFPOSX1 \RF_reg[22][13]  ( .D(n2784), .CLK(clk), .Q(\RF[22][13] ) );
  DFFPOSX1 \RF_reg[22][12]  ( .D(n2783), .CLK(clk), .Q(\RF[22][12] ) );
  DFFPOSX1 \RF_reg[22][11]  ( .D(n2782), .CLK(clk), .Q(\RF[22][11] ) );
  DFFPOSX1 \RF_reg[22][10]  ( .D(n2781), .CLK(clk), .Q(\RF[22][10] ) );
  DFFPOSX1 \RF_reg[22][9]  ( .D(n2780), .CLK(clk), .Q(\RF[22][9] ) );
  DFFPOSX1 \RF_reg[22][8]  ( .D(n2779), .CLK(clk), .Q(\RF[22][8] ) );
  DFFPOSX1 \RF_reg[22][7]  ( .D(n2778), .CLK(clk), .Q(\RF[22][7] ) );
  DFFPOSX1 \RF_reg[22][6]  ( .D(n2777), .CLK(clk), .Q(\RF[22][6] ) );
  DFFPOSX1 \RF_reg[22][5]  ( .D(n2776), .CLK(clk), .Q(\RF[22][5] ) );
  DFFPOSX1 \RF_reg[22][4]  ( .D(n2775), .CLK(clk), .Q(\RF[22][4] ) );
  DFFPOSX1 \RF_reg[22][3]  ( .D(n2774), .CLK(clk), .Q(\RF[22][3] ) );
  DFFPOSX1 \RF_reg[22][2]  ( .D(n2773), .CLK(clk), .Q(\RF[22][2] ) );
  DFFPOSX1 \RF_reg[22][1]  ( .D(n2772), .CLK(clk), .Q(\RF[22][1] ) );
  DFFPOSX1 \RF_reg[22][0]  ( .D(n2771), .CLK(clk), .Q(\RF[22][0] ) );
  DFFPOSX1 \RF_reg[23][63]  ( .D(n2770), .CLK(clk), .Q(\RF[23][63] ) );
  DFFPOSX1 \RF_reg[23][62]  ( .D(n2769), .CLK(clk), .Q(\RF[23][62] ) );
  DFFPOSX1 \RF_reg[23][61]  ( .D(n2768), .CLK(clk), .Q(\RF[23][61] ) );
  DFFPOSX1 \RF_reg[23][60]  ( .D(n2767), .CLK(clk), .Q(\RF[23][60] ) );
  DFFPOSX1 \RF_reg[23][59]  ( .D(n2766), .CLK(clk), .Q(\RF[23][59] ) );
  DFFPOSX1 \RF_reg[23][58]  ( .D(n2765), .CLK(clk), .Q(\RF[23][58] ) );
  DFFPOSX1 \RF_reg[23][57]  ( .D(n2764), .CLK(clk), .Q(\RF[23][57] ) );
  DFFPOSX1 \RF_reg[23][56]  ( .D(n2763), .CLK(clk), .Q(\RF[23][56] ) );
  DFFPOSX1 \RF_reg[23][55]  ( .D(n2762), .CLK(clk), .Q(\RF[23][55] ) );
  DFFPOSX1 \RF_reg[23][54]  ( .D(n2761), .CLK(clk), .Q(\RF[23][54] ) );
  DFFPOSX1 \RF_reg[23][53]  ( .D(n2760), .CLK(clk), .Q(\RF[23][53] ) );
  DFFPOSX1 \RF_reg[23][52]  ( .D(n2759), .CLK(clk), .Q(\RF[23][52] ) );
  DFFPOSX1 \RF_reg[23][51]  ( .D(n2758), .CLK(clk), .Q(\RF[23][51] ) );
  DFFPOSX1 \RF_reg[23][50]  ( .D(n2757), .CLK(clk), .Q(\RF[23][50] ) );
  DFFPOSX1 \RF_reg[23][49]  ( .D(n2756), .CLK(clk), .Q(\RF[23][49] ) );
  DFFPOSX1 \RF_reg[23][48]  ( .D(n2755), .CLK(clk), .Q(\RF[23][48] ) );
  DFFPOSX1 \RF_reg[23][47]  ( .D(n2754), .CLK(clk), .Q(\RF[23][47] ) );
  DFFPOSX1 \RF_reg[23][46]  ( .D(n2753), .CLK(clk), .Q(\RF[23][46] ) );
  DFFPOSX1 \RF_reg[23][45]  ( .D(n2752), .CLK(clk), .Q(\RF[23][45] ) );
  DFFPOSX1 \RF_reg[23][44]  ( .D(n2751), .CLK(clk), .Q(\RF[23][44] ) );
  DFFPOSX1 \RF_reg[23][43]  ( .D(n2750), .CLK(clk), .Q(\RF[23][43] ) );
  DFFPOSX1 \RF_reg[23][42]  ( .D(n2749), .CLK(clk), .Q(\RF[23][42] ) );
  DFFPOSX1 \RF_reg[23][41]  ( .D(n2748), .CLK(clk), .Q(\RF[23][41] ) );
  DFFPOSX1 \RF_reg[23][40]  ( .D(n2747), .CLK(clk), .Q(\RF[23][40] ) );
  DFFPOSX1 \RF_reg[23][39]  ( .D(n2746), .CLK(clk), .Q(\RF[23][39] ) );
  DFFPOSX1 \RF_reg[23][38]  ( .D(n2745), .CLK(clk), .Q(\RF[23][38] ) );
  DFFPOSX1 \RF_reg[23][37]  ( .D(n2744), .CLK(clk), .Q(\RF[23][37] ) );
  DFFPOSX1 \RF_reg[23][36]  ( .D(n2743), .CLK(clk), .Q(\RF[23][36] ) );
  DFFPOSX1 \RF_reg[23][35]  ( .D(n2742), .CLK(clk), .Q(\RF[23][35] ) );
  DFFPOSX1 \RF_reg[23][34]  ( .D(n2741), .CLK(clk), .Q(\RF[23][34] ) );
  DFFPOSX1 \RF_reg[23][33]  ( .D(n2740), .CLK(clk), .Q(\RF[23][33] ) );
  DFFPOSX1 \RF_reg[23][32]  ( .D(n2739), .CLK(clk), .Q(\RF[23][32] ) );
  DFFPOSX1 \RF_reg[23][31]  ( .D(n2738), .CLK(clk), .Q(\RF[23][31] ) );
  DFFPOSX1 \RF_reg[23][30]  ( .D(n2737), .CLK(clk), .Q(\RF[23][30] ) );
  DFFPOSX1 \RF_reg[23][29]  ( .D(n2736), .CLK(clk), .Q(\RF[23][29] ) );
  DFFPOSX1 \RF_reg[23][28]  ( .D(n2735), .CLK(clk), .Q(\RF[23][28] ) );
  DFFPOSX1 \RF_reg[23][27]  ( .D(n2734), .CLK(clk), .Q(\RF[23][27] ) );
  DFFPOSX1 \RF_reg[23][26]  ( .D(n2733), .CLK(clk), .Q(\RF[23][26] ) );
  DFFPOSX1 \RF_reg[23][25]  ( .D(n2732), .CLK(clk), .Q(\RF[23][25] ) );
  DFFPOSX1 \RF_reg[23][24]  ( .D(n2731), .CLK(clk), .Q(\RF[23][24] ) );
  DFFPOSX1 \RF_reg[23][23]  ( .D(n2730), .CLK(clk), .Q(\RF[23][23] ) );
  DFFPOSX1 \RF_reg[23][22]  ( .D(n2729), .CLK(clk), .Q(\RF[23][22] ) );
  DFFPOSX1 \RF_reg[23][21]  ( .D(n2728), .CLK(clk), .Q(\RF[23][21] ) );
  DFFPOSX1 \RF_reg[23][20]  ( .D(n2727), .CLK(clk), .Q(\RF[23][20] ) );
  DFFPOSX1 \RF_reg[23][19]  ( .D(n2726), .CLK(clk), .Q(\RF[23][19] ) );
  DFFPOSX1 \RF_reg[23][18]  ( .D(n2725), .CLK(clk), .Q(\RF[23][18] ) );
  DFFPOSX1 \RF_reg[23][17]  ( .D(n2724), .CLK(clk), .Q(\RF[23][17] ) );
  DFFPOSX1 \RF_reg[23][16]  ( .D(n2723), .CLK(clk), .Q(\RF[23][16] ) );
  DFFPOSX1 \RF_reg[23][15]  ( .D(n2722), .CLK(clk), .Q(\RF[23][15] ) );
  DFFPOSX1 \RF_reg[23][14]  ( .D(n2721), .CLK(clk), .Q(\RF[23][14] ) );
  DFFPOSX1 \RF_reg[23][13]  ( .D(n2720), .CLK(clk), .Q(\RF[23][13] ) );
  DFFPOSX1 \RF_reg[23][12]  ( .D(n2719), .CLK(clk), .Q(\RF[23][12] ) );
  DFFPOSX1 \RF_reg[23][11]  ( .D(n2718), .CLK(clk), .Q(\RF[23][11] ) );
  DFFPOSX1 \RF_reg[23][10]  ( .D(n2717), .CLK(clk), .Q(\RF[23][10] ) );
  DFFPOSX1 \RF_reg[23][9]  ( .D(n2716), .CLK(clk), .Q(\RF[23][9] ) );
  DFFPOSX1 \RF_reg[23][8]  ( .D(n2715), .CLK(clk), .Q(\RF[23][8] ) );
  DFFPOSX1 \RF_reg[23][7]  ( .D(n2714), .CLK(clk), .Q(\RF[23][7] ) );
  DFFPOSX1 \RF_reg[23][6]  ( .D(n2713), .CLK(clk), .Q(\RF[23][6] ) );
  DFFPOSX1 \RF_reg[23][5]  ( .D(n2712), .CLK(clk), .Q(\RF[23][5] ) );
  DFFPOSX1 \RF_reg[23][4]  ( .D(n2711), .CLK(clk), .Q(\RF[23][4] ) );
  DFFPOSX1 \RF_reg[23][3]  ( .D(n2710), .CLK(clk), .Q(\RF[23][3] ) );
  DFFPOSX1 \RF_reg[23][2]  ( .D(n2709), .CLK(clk), .Q(\RF[23][2] ) );
  DFFPOSX1 \RF_reg[23][1]  ( .D(n2708), .CLK(clk), .Q(\RF[23][1] ) );
  DFFPOSX1 \RF_reg[23][0]  ( .D(n2707), .CLK(clk), .Q(\RF[23][0] ) );
  DFFPOSX1 \RF_reg[24][63]  ( .D(n2706), .CLK(clk), .Q(\RF[24][63] ) );
  DFFPOSX1 \RF_reg[24][62]  ( .D(n2705), .CLK(clk), .Q(\RF[24][62] ) );
  DFFPOSX1 \RF_reg[24][61]  ( .D(n2704), .CLK(clk), .Q(\RF[24][61] ) );
  DFFPOSX1 \RF_reg[24][60]  ( .D(n2703), .CLK(clk), .Q(\RF[24][60] ) );
  DFFPOSX1 \RF_reg[24][59]  ( .D(n2702), .CLK(clk), .Q(\RF[24][59] ) );
  DFFPOSX1 \RF_reg[24][58]  ( .D(n2701), .CLK(clk), .Q(\RF[24][58] ) );
  DFFPOSX1 \RF_reg[24][57]  ( .D(n2700), .CLK(clk), .Q(\RF[24][57] ) );
  DFFPOSX1 \RF_reg[24][56]  ( .D(n2699), .CLK(clk), .Q(\RF[24][56] ) );
  DFFPOSX1 \RF_reg[24][55]  ( .D(n2698), .CLK(clk), .Q(\RF[24][55] ) );
  DFFPOSX1 \RF_reg[24][54]  ( .D(n2697), .CLK(clk), .Q(\RF[24][54] ) );
  DFFPOSX1 \RF_reg[24][53]  ( .D(n2696), .CLK(clk), .Q(\RF[24][53] ) );
  DFFPOSX1 \RF_reg[24][52]  ( .D(n2695), .CLK(clk), .Q(\RF[24][52] ) );
  DFFPOSX1 \RF_reg[24][51]  ( .D(n2694), .CLK(clk), .Q(\RF[24][51] ) );
  DFFPOSX1 \RF_reg[24][50]  ( .D(n2693), .CLK(clk), .Q(\RF[24][50] ) );
  DFFPOSX1 \RF_reg[24][49]  ( .D(n2692), .CLK(clk), .Q(\RF[24][49] ) );
  DFFPOSX1 \RF_reg[24][48]  ( .D(n2691), .CLK(clk), .Q(\RF[24][48] ) );
  DFFPOSX1 \RF_reg[24][47]  ( .D(n2690), .CLK(clk), .Q(\RF[24][47] ) );
  DFFPOSX1 \RF_reg[24][46]  ( .D(n2689), .CLK(clk), .Q(\RF[24][46] ) );
  DFFPOSX1 \RF_reg[24][45]  ( .D(n2688), .CLK(clk), .Q(\RF[24][45] ) );
  DFFPOSX1 \RF_reg[24][44]  ( .D(n2687), .CLK(clk), .Q(\RF[24][44] ) );
  DFFPOSX1 \RF_reg[24][43]  ( .D(n2686), .CLK(clk), .Q(\RF[24][43] ) );
  DFFPOSX1 \RF_reg[24][42]  ( .D(n2685), .CLK(clk), .Q(\RF[24][42] ) );
  DFFPOSX1 \RF_reg[24][41]  ( .D(n2684), .CLK(clk), .Q(\RF[24][41] ) );
  DFFPOSX1 \RF_reg[24][40]  ( .D(n2683), .CLK(clk), .Q(\RF[24][40] ) );
  DFFPOSX1 \RF_reg[24][39]  ( .D(n2682), .CLK(clk), .Q(\RF[24][39] ) );
  DFFPOSX1 \RF_reg[24][38]  ( .D(n2681), .CLK(clk), .Q(\RF[24][38] ) );
  DFFPOSX1 \RF_reg[24][37]  ( .D(n2680), .CLK(clk), .Q(\RF[24][37] ) );
  DFFPOSX1 \RF_reg[24][36]  ( .D(n2679), .CLK(clk), .Q(\RF[24][36] ) );
  DFFPOSX1 \RF_reg[24][35]  ( .D(n2678), .CLK(clk), .Q(\RF[24][35] ) );
  DFFPOSX1 \RF_reg[24][34]  ( .D(n2677), .CLK(clk), .Q(\RF[24][34] ) );
  DFFPOSX1 \RF_reg[24][33]  ( .D(n2676), .CLK(clk), .Q(\RF[24][33] ) );
  DFFPOSX1 \RF_reg[24][32]  ( .D(n2675), .CLK(clk), .Q(\RF[24][32] ) );
  DFFPOSX1 \RF_reg[24][31]  ( .D(n2674), .CLK(clk), .Q(\RF[24][31] ) );
  DFFPOSX1 \RF_reg[24][30]  ( .D(n2673), .CLK(clk), .Q(\RF[24][30] ) );
  DFFPOSX1 \RF_reg[24][29]  ( .D(n2672), .CLK(clk), .Q(\RF[24][29] ) );
  DFFPOSX1 \RF_reg[24][28]  ( .D(n2671), .CLK(clk), .Q(\RF[24][28] ) );
  DFFPOSX1 \RF_reg[24][27]  ( .D(n2670), .CLK(clk), .Q(\RF[24][27] ) );
  DFFPOSX1 \RF_reg[24][26]  ( .D(n2669), .CLK(clk), .Q(\RF[24][26] ) );
  DFFPOSX1 \RF_reg[24][25]  ( .D(n2668), .CLK(clk), .Q(\RF[24][25] ) );
  DFFPOSX1 \RF_reg[24][24]  ( .D(n2667), .CLK(clk), .Q(\RF[24][24] ) );
  DFFPOSX1 \RF_reg[24][23]  ( .D(n2666), .CLK(clk), .Q(\RF[24][23] ) );
  DFFPOSX1 \RF_reg[24][22]  ( .D(n2665), .CLK(clk), .Q(\RF[24][22] ) );
  DFFPOSX1 \RF_reg[24][21]  ( .D(n2664), .CLK(clk), .Q(\RF[24][21] ) );
  DFFPOSX1 \RF_reg[24][20]  ( .D(n2663), .CLK(clk), .Q(\RF[24][20] ) );
  DFFPOSX1 \RF_reg[24][19]  ( .D(n2662), .CLK(clk), .Q(\RF[24][19] ) );
  DFFPOSX1 \RF_reg[24][18]  ( .D(n2661), .CLK(clk), .Q(\RF[24][18] ) );
  DFFPOSX1 \RF_reg[24][17]  ( .D(n2660), .CLK(clk), .Q(\RF[24][17] ) );
  DFFPOSX1 \RF_reg[24][16]  ( .D(n2659), .CLK(clk), .Q(\RF[24][16] ) );
  DFFPOSX1 \RF_reg[24][15]  ( .D(n2658), .CLK(clk), .Q(\RF[24][15] ) );
  DFFPOSX1 \RF_reg[24][14]  ( .D(n2657), .CLK(clk), .Q(\RF[24][14] ) );
  DFFPOSX1 \RF_reg[24][13]  ( .D(n2656), .CLK(clk), .Q(\RF[24][13] ) );
  DFFPOSX1 \RF_reg[24][12]  ( .D(n2655), .CLK(clk), .Q(\RF[24][12] ) );
  DFFPOSX1 \RF_reg[24][11]  ( .D(n2654), .CLK(clk), .Q(\RF[24][11] ) );
  DFFPOSX1 \RF_reg[24][10]  ( .D(n2653), .CLK(clk), .Q(\RF[24][10] ) );
  DFFPOSX1 \RF_reg[24][9]  ( .D(n2652), .CLK(clk), .Q(\RF[24][9] ) );
  DFFPOSX1 \RF_reg[24][8]  ( .D(n2651), .CLK(clk), .Q(\RF[24][8] ) );
  DFFPOSX1 \RF_reg[24][7]  ( .D(n2650), .CLK(clk), .Q(\RF[24][7] ) );
  DFFPOSX1 \RF_reg[24][6]  ( .D(n2649), .CLK(clk), .Q(\RF[24][6] ) );
  DFFPOSX1 \RF_reg[24][5]  ( .D(n2648), .CLK(clk), .Q(\RF[24][5] ) );
  DFFPOSX1 \RF_reg[24][4]  ( .D(n2647), .CLK(clk), .Q(\RF[24][4] ) );
  DFFPOSX1 \RF_reg[24][3]  ( .D(n2646), .CLK(clk), .Q(\RF[24][3] ) );
  DFFPOSX1 \RF_reg[24][2]  ( .D(n2645), .CLK(clk), .Q(\RF[24][2] ) );
  DFFPOSX1 \RF_reg[24][1]  ( .D(n2644), .CLK(clk), .Q(\RF[24][1] ) );
  DFFPOSX1 \RF_reg[24][0]  ( .D(n2643), .CLK(clk), .Q(\RF[24][0] ) );
  DFFPOSX1 \RF_reg[25][63]  ( .D(n2642), .CLK(clk), .Q(\RF[25][63] ) );
  DFFPOSX1 \RF_reg[25][62]  ( .D(n2641), .CLK(clk), .Q(\RF[25][62] ) );
  DFFPOSX1 \RF_reg[25][61]  ( .D(n2640), .CLK(clk), .Q(\RF[25][61] ) );
  DFFPOSX1 \RF_reg[25][60]  ( .D(n2639), .CLK(clk), .Q(\RF[25][60] ) );
  DFFPOSX1 \RF_reg[25][59]  ( .D(n2638), .CLK(clk), .Q(\RF[25][59] ) );
  DFFPOSX1 \RF_reg[25][58]  ( .D(n2637), .CLK(clk), .Q(\RF[25][58] ) );
  DFFPOSX1 \RF_reg[25][57]  ( .D(n2636), .CLK(clk), .Q(\RF[25][57] ) );
  DFFPOSX1 \RF_reg[25][56]  ( .D(n2635), .CLK(clk), .Q(\RF[25][56] ) );
  DFFPOSX1 \RF_reg[25][55]  ( .D(n2634), .CLK(clk), .Q(\RF[25][55] ) );
  DFFPOSX1 \RF_reg[25][54]  ( .D(n2633), .CLK(clk), .Q(\RF[25][54] ) );
  DFFPOSX1 \RF_reg[25][53]  ( .D(n2632), .CLK(clk), .Q(\RF[25][53] ) );
  DFFPOSX1 \RF_reg[25][52]  ( .D(n2631), .CLK(clk), .Q(\RF[25][52] ) );
  DFFPOSX1 \RF_reg[25][51]  ( .D(n2630), .CLK(clk), .Q(\RF[25][51] ) );
  DFFPOSX1 \RF_reg[25][50]  ( .D(n2629), .CLK(clk), .Q(\RF[25][50] ) );
  DFFPOSX1 \RF_reg[25][49]  ( .D(n2628), .CLK(clk), .Q(\RF[25][49] ) );
  DFFPOSX1 \RF_reg[25][48]  ( .D(n2627), .CLK(clk), .Q(\RF[25][48] ) );
  DFFPOSX1 \RF_reg[25][47]  ( .D(n2626), .CLK(clk), .Q(\RF[25][47] ) );
  DFFPOSX1 \RF_reg[25][46]  ( .D(n2625), .CLK(clk), .Q(\RF[25][46] ) );
  DFFPOSX1 \RF_reg[25][45]  ( .D(n2624), .CLK(clk), .Q(\RF[25][45] ) );
  DFFPOSX1 \RF_reg[25][44]  ( .D(n2623), .CLK(clk), .Q(\RF[25][44] ) );
  DFFPOSX1 \RF_reg[25][43]  ( .D(n2622), .CLK(clk), .Q(\RF[25][43] ) );
  DFFPOSX1 \RF_reg[25][42]  ( .D(n2621), .CLK(clk), .Q(\RF[25][42] ) );
  DFFPOSX1 \RF_reg[25][41]  ( .D(n2620), .CLK(clk), .Q(\RF[25][41] ) );
  DFFPOSX1 \RF_reg[25][40]  ( .D(n2619), .CLK(clk), .Q(\RF[25][40] ) );
  DFFPOSX1 \RF_reg[25][39]  ( .D(n2618), .CLK(clk), .Q(\RF[25][39] ) );
  DFFPOSX1 \RF_reg[25][38]  ( .D(n2617), .CLK(clk), .Q(\RF[25][38] ) );
  DFFPOSX1 \RF_reg[25][37]  ( .D(n2616), .CLK(clk), .Q(\RF[25][37] ) );
  DFFPOSX1 \RF_reg[25][36]  ( .D(n2615), .CLK(clk), .Q(\RF[25][36] ) );
  DFFPOSX1 \RF_reg[25][35]  ( .D(n2614), .CLK(clk), .Q(\RF[25][35] ) );
  DFFPOSX1 \RF_reg[25][34]  ( .D(n2613), .CLK(clk), .Q(\RF[25][34] ) );
  DFFPOSX1 \RF_reg[25][33]  ( .D(n2612), .CLK(clk), .Q(\RF[25][33] ) );
  DFFPOSX1 \RF_reg[25][32]  ( .D(n2611), .CLK(clk), .Q(\RF[25][32] ) );
  DFFPOSX1 \RF_reg[25][31]  ( .D(n2610), .CLK(clk), .Q(\RF[25][31] ) );
  DFFPOSX1 \RF_reg[25][30]  ( .D(n2609), .CLK(clk), .Q(\RF[25][30] ) );
  DFFPOSX1 \RF_reg[25][29]  ( .D(n2608), .CLK(clk), .Q(\RF[25][29] ) );
  DFFPOSX1 \RF_reg[25][28]  ( .D(n2607), .CLK(clk), .Q(\RF[25][28] ) );
  DFFPOSX1 \RF_reg[25][27]  ( .D(n2606), .CLK(clk), .Q(\RF[25][27] ) );
  DFFPOSX1 \RF_reg[25][26]  ( .D(n2605), .CLK(clk), .Q(\RF[25][26] ) );
  DFFPOSX1 \RF_reg[25][25]  ( .D(n2604), .CLK(clk), .Q(\RF[25][25] ) );
  DFFPOSX1 \RF_reg[25][24]  ( .D(n2603), .CLK(clk), .Q(\RF[25][24] ) );
  DFFPOSX1 \RF_reg[25][23]  ( .D(n2602), .CLK(clk), .Q(\RF[25][23] ) );
  DFFPOSX1 \RF_reg[25][22]  ( .D(n2601), .CLK(clk), .Q(\RF[25][22] ) );
  DFFPOSX1 \RF_reg[25][21]  ( .D(n2600), .CLK(clk), .Q(\RF[25][21] ) );
  DFFPOSX1 \RF_reg[25][20]  ( .D(n2599), .CLK(clk), .Q(\RF[25][20] ) );
  DFFPOSX1 \RF_reg[25][19]  ( .D(n2598), .CLK(clk), .Q(\RF[25][19] ) );
  DFFPOSX1 \RF_reg[25][18]  ( .D(n2597), .CLK(clk), .Q(\RF[25][18] ) );
  DFFPOSX1 \RF_reg[25][17]  ( .D(n2596), .CLK(clk), .Q(\RF[25][17] ) );
  DFFPOSX1 \RF_reg[25][16]  ( .D(n2595), .CLK(clk), .Q(\RF[25][16] ) );
  DFFPOSX1 \RF_reg[25][15]  ( .D(n2594), .CLK(clk), .Q(\RF[25][15] ) );
  DFFPOSX1 \RF_reg[25][14]  ( .D(n2593), .CLK(clk), .Q(\RF[25][14] ) );
  DFFPOSX1 \RF_reg[25][13]  ( .D(n2592), .CLK(clk), .Q(\RF[25][13] ) );
  DFFPOSX1 \RF_reg[25][12]  ( .D(n2591), .CLK(clk), .Q(\RF[25][12] ) );
  DFFPOSX1 \RF_reg[25][11]  ( .D(n2590), .CLK(clk), .Q(\RF[25][11] ) );
  DFFPOSX1 \RF_reg[25][10]  ( .D(n2589), .CLK(clk), .Q(\RF[25][10] ) );
  DFFPOSX1 \RF_reg[25][9]  ( .D(n2588), .CLK(clk), .Q(\RF[25][9] ) );
  DFFPOSX1 \RF_reg[25][8]  ( .D(n2587), .CLK(clk), .Q(\RF[25][8] ) );
  DFFPOSX1 \RF_reg[25][7]  ( .D(n2586), .CLK(clk), .Q(\RF[25][7] ) );
  DFFPOSX1 \RF_reg[25][6]  ( .D(n2585), .CLK(clk), .Q(\RF[25][6] ) );
  DFFPOSX1 \RF_reg[25][5]  ( .D(n2584), .CLK(clk), .Q(\RF[25][5] ) );
  DFFPOSX1 \RF_reg[25][4]  ( .D(n2583), .CLK(clk), .Q(\RF[25][4] ) );
  DFFPOSX1 \RF_reg[25][3]  ( .D(n2582), .CLK(clk), .Q(\RF[25][3] ) );
  DFFPOSX1 \RF_reg[25][2]  ( .D(n2581), .CLK(clk), .Q(\RF[25][2] ) );
  DFFPOSX1 \RF_reg[25][1]  ( .D(n2580), .CLK(clk), .Q(\RF[25][1] ) );
  DFFPOSX1 \RF_reg[25][0]  ( .D(n2579), .CLK(clk), .Q(\RF[25][0] ) );
  DFFPOSX1 \RF_reg[26][63]  ( .D(n2578), .CLK(clk), .Q(\RF[26][63] ) );
  DFFPOSX1 \RF_reg[26][62]  ( .D(n2577), .CLK(clk), .Q(\RF[26][62] ) );
  DFFPOSX1 \RF_reg[26][61]  ( .D(n2576), .CLK(clk), .Q(\RF[26][61] ) );
  DFFPOSX1 \RF_reg[26][60]  ( .D(n2575), .CLK(clk), .Q(\RF[26][60] ) );
  DFFPOSX1 \RF_reg[26][59]  ( .D(n2574), .CLK(clk), .Q(\RF[26][59] ) );
  DFFPOSX1 \RF_reg[26][58]  ( .D(n2573), .CLK(clk), .Q(\RF[26][58] ) );
  DFFPOSX1 \RF_reg[26][57]  ( .D(n2572), .CLK(clk), .Q(\RF[26][57] ) );
  DFFPOSX1 \RF_reg[26][56]  ( .D(n2571), .CLK(clk), .Q(\RF[26][56] ) );
  DFFPOSX1 \RF_reg[26][55]  ( .D(n2570), .CLK(clk), .Q(\RF[26][55] ) );
  DFFPOSX1 \RF_reg[26][54]  ( .D(n2569), .CLK(clk), .Q(\RF[26][54] ) );
  DFFPOSX1 \RF_reg[26][53]  ( .D(n2568), .CLK(clk), .Q(\RF[26][53] ) );
  DFFPOSX1 \RF_reg[26][52]  ( .D(n2567), .CLK(clk), .Q(\RF[26][52] ) );
  DFFPOSX1 \RF_reg[26][51]  ( .D(n2566), .CLK(clk), .Q(\RF[26][51] ) );
  DFFPOSX1 \RF_reg[26][50]  ( .D(n2565), .CLK(clk), .Q(\RF[26][50] ) );
  DFFPOSX1 \RF_reg[26][49]  ( .D(n2564), .CLK(clk), .Q(\RF[26][49] ) );
  DFFPOSX1 \RF_reg[26][48]  ( .D(n2563), .CLK(clk), .Q(\RF[26][48] ) );
  DFFPOSX1 \RF_reg[26][47]  ( .D(n2562), .CLK(clk), .Q(\RF[26][47] ) );
  DFFPOSX1 \RF_reg[26][46]  ( .D(n2561), .CLK(clk), .Q(\RF[26][46] ) );
  DFFPOSX1 \RF_reg[26][45]  ( .D(n2560), .CLK(clk), .Q(\RF[26][45] ) );
  DFFPOSX1 \RF_reg[26][44]  ( .D(n2559), .CLK(clk), .Q(\RF[26][44] ) );
  DFFPOSX1 \RF_reg[26][43]  ( .D(n2558), .CLK(clk), .Q(\RF[26][43] ) );
  DFFPOSX1 \RF_reg[26][42]  ( .D(n2557), .CLK(clk), .Q(\RF[26][42] ) );
  DFFPOSX1 \RF_reg[26][41]  ( .D(n2556), .CLK(clk), .Q(\RF[26][41] ) );
  DFFPOSX1 \RF_reg[26][40]  ( .D(n2555), .CLK(clk), .Q(\RF[26][40] ) );
  DFFPOSX1 \RF_reg[26][39]  ( .D(n2554), .CLK(clk), .Q(\RF[26][39] ) );
  DFFPOSX1 \RF_reg[26][38]  ( .D(n2553), .CLK(clk), .Q(\RF[26][38] ) );
  DFFPOSX1 \RF_reg[26][37]  ( .D(n2552), .CLK(clk), .Q(\RF[26][37] ) );
  DFFPOSX1 \RF_reg[26][36]  ( .D(n2551), .CLK(clk), .Q(\RF[26][36] ) );
  DFFPOSX1 \RF_reg[26][35]  ( .D(n2550), .CLK(clk), .Q(\RF[26][35] ) );
  DFFPOSX1 \RF_reg[26][34]  ( .D(n2549), .CLK(clk), .Q(\RF[26][34] ) );
  DFFPOSX1 \RF_reg[26][33]  ( .D(n2548), .CLK(clk), .Q(\RF[26][33] ) );
  DFFPOSX1 \RF_reg[26][32]  ( .D(n2547), .CLK(clk), .Q(\RF[26][32] ) );
  DFFPOSX1 \RF_reg[26][31]  ( .D(n2546), .CLK(clk), .Q(\RF[26][31] ) );
  DFFPOSX1 \RF_reg[26][30]  ( .D(n2545), .CLK(clk), .Q(\RF[26][30] ) );
  DFFPOSX1 \RF_reg[26][29]  ( .D(n2544), .CLK(clk), .Q(\RF[26][29] ) );
  DFFPOSX1 \RF_reg[26][28]  ( .D(n2543), .CLK(clk), .Q(\RF[26][28] ) );
  DFFPOSX1 \RF_reg[26][27]  ( .D(n2542), .CLK(clk), .Q(\RF[26][27] ) );
  DFFPOSX1 \RF_reg[26][26]  ( .D(n2541), .CLK(clk), .Q(\RF[26][26] ) );
  DFFPOSX1 \RF_reg[26][25]  ( .D(n2540), .CLK(clk), .Q(\RF[26][25] ) );
  DFFPOSX1 \RF_reg[26][24]  ( .D(n2539), .CLK(clk), .Q(\RF[26][24] ) );
  DFFPOSX1 \RF_reg[26][23]  ( .D(n2538), .CLK(clk), .Q(\RF[26][23] ) );
  DFFPOSX1 \RF_reg[26][22]  ( .D(n2537), .CLK(clk), .Q(\RF[26][22] ) );
  DFFPOSX1 \RF_reg[26][21]  ( .D(n2536), .CLK(clk), .Q(\RF[26][21] ) );
  DFFPOSX1 \RF_reg[26][20]  ( .D(n2535), .CLK(clk), .Q(\RF[26][20] ) );
  DFFPOSX1 \RF_reg[26][19]  ( .D(n2534), .CLK(clk), .Q(\RF[26][19] ) );
  DFFPOSX1 \RF_reg[26][18]  ( .D(n2533), .CLK(clk), .Q(\RF[26][18] ) );
  DFFPOSX1 \RF_reg[26][17]  ( .D(n2532), .CLK(clk), .Q(\RF[26][17] ) );
  DFFPOSX1 \RF_reg[26][16]  ( .D(n2531), .CLK(clk), .Q(\RF[26][16] ) );
  DFFPOSX1 \RF_reg[26][15]  ( .D(n2530), .CLK(clk), .Q(\RF[26][15] ) );
  DFFPOSX1 \RF_reg[26][14]  ( .D(n2529), .CLK(clk), .Q(\RF[26][14] ) );
  DFFPOSX1 \RF_reg[26][13]  ( .D(n2528), .CLK(clk), .Q(\RF[26][13] ) );
  DFFPOSX1 \RF_reg[26][12]  ( .D(n2527), .CLK(clk), .Q(\RF[26][12] ) );
  DFFPOSX1 \RF_reg[26][11]  ( .D(n2526), .CLK(clk), .Q(\RF[26][11] ) );
  DFFPOSX1 \RF_reg[26][10]  ( .D(n2525), .CLK(clk), .Q(\RF[26][10] ) );
  DFFPOSX1 \RF_reg[26][9]  ( .D(n2524), .CLK(clk), .Q(\RF[26][9] ) );
  DFFPOSX1 \RF_reg[26][8]  ( .D(n2523), .CLK(clk), .Q(\RF[26][8] ) );
  DFFPOSX1 \RF_reg[26][7]  ( .D(n2522), .CLK(clk), .Q(\RF[26][7] ) );
  DFFPOSX1 \RF_reg[26][6]  ( .D(n2521), .CLK(clk), .Q(\RF[26][6] ) );
  DFFPOSX1 \RF_reg[26][5]  ( .D(n2520), .CLK(clk), .Q(\RF[26][5] ) );
  DFFPOSX1 \RF_reg[26][4]  ( .D(n2519), .CLK(clk), .Q(\RF[26][4] ) );
  DFFPOSX1 \RF_reg[26][3]  ( .D(n2518), .CLK(clk), .Q(\RF[26][3] ) );
  DFFPOSX1 \RF_reg[26][2]  ( .D(n2517), .CLK(clk), .Q(\RF[26][2] ) );
  DFFPOSX1 \RF_reg[26][1]  ( .D(n2516), .CLK(clk), .Q(\RF[26][1] ) );
  DFFPOSX1 \RF_reg[26][0]  ( .D(n2515), .CLK(clk), .Q(\RF[26][0] ) );
  DFFPOSX1 \RF_reg[27][63]  ( .D(n2514), .CLK(clk), .Q(\RF[27][63] ) );
  DFFPOSX1 \RF_reg[27][62]  ( .D(n2513), .CLK(clk), .Q(\RF[27][62] ) );
  DFFPOSX1 \RF_reg[27][61]  ( .D(n2512), .CLK(clk), .Q(\RF[27][61] ) );
  DFFPOSX1 \RF_reg[27][60]  ( .D(n2511), .CLK(clk), .Q(\RF[27][60] ) );
  DFFPOSX1 \RF_reg[27][59]  ( .D(n2510), .CLK(clk), .Q(\RF[27][59] ) );
  DFFPOSX1 \RF_reg[27][58]  ( .D(n2509), .CLK(clk), .Q(\RF[27][58] ) );
  DFFPOSX1 \RF_reg[27][57]  ( .D(n2508), .CLK(clk), .Q(\RF[27][57] ) );
  DFFPOSX1 \RF_reg[27][56]  ( .D(n2507), .CLK(clk), .Q(\RF[27][56] ) );
  DFFPOSX1 \RF_reg[27][55]  ( .D(n2506), .CLK(clk), .Q(\RF[27][55] ) );
  DFFPOSX1 \RF_reg[27][54]  ( .D(n2505), .CLK(clk), .Q(\RF[27][54] ) );
  DFFPOSX1 \RF_reg[27][53]  ( .D(n2504), .CLK(clk), .Q(\RF[27][53] ) );
  DFFPOSX1 \RF_reg[27][52]  ( .D(n2503), .CLK(clk), .Q(\RF[27][52] ) );
  DFFPOSX1 \RF_reg[27][51]  ( .D(n2502), .CLK(clk), .Q(\RF[27][51] ) );
  DFFPOSX1 \RF_reg[27][50]  ( .D(n2501), .CLK(clk), .Q(\RF[27][50] ) );
  DFFPOSX1 \RF_reg[27][49]  ( .D(n2500), .CLK(clk), .Q(\RF[27][49] ) );
  DFFPOSX1 \RF_reg[27][48]  ( .D(n2499), .CLK(clk), .Q(\RF[27][48] ) );
  DFFPOSX1 \RF_reg[27][47]  ( .D(n2498), .CLK(clk), .Q(\RF[27][47] ) );
  DFFPOSX1 \RF_reg[27][46]  ( .D(n2497), .CLK(clk), .Q(\RF[27][46] ) );
  DFFPOSX1 \RF_reg[27][45]  ( .D(n2496), .CLK(clk), .Q(\RF[27][45] ) );
  DFFPOSX1 \RF_reg[27][44]  ( .D(n2495), .CLK(clk), .Q(\RF[27][44] ) );
  DFFPOSX1 \RF_reg[27][43]  ( .D(n2494), .CLK(clk), .Q(\RF[27][43] ) );
  DFFPOSX1 \RF_reg[27][42]  ( .D(n2493), .CLK(clk), .Q(\RF[27][42] ) );
  DFFPOSX1 \RF_reg[27][41]  ( .D(n2492), .CLK(clk), .Q(\RF[27][41] ) );
  DFFPOSX1 \RF_reg[27][40]  ( .D(n2491), .CLK(clk), .Q(\RF[27][40] ) );
  DFFPOSX1 \RF_reg[27][39]  ( .D(n2490), .CLK(clk), .Q(\RF[27][39] ) );
  DFFPOSX1 \RF_reg[27][38]  ( .D(n2489), .CLK(clk), .Q(\RF[27][38] ) );
  DFFPOSX1 \RF_reg[27][37]  ( .D(n2488), .CLK(clk), .Q(\RF[27][37] ) );
  DFFPOSX1 \RF_reg[27][36]  ( .D(n2487), .CLK(clk), .Q(\RF[27][36] ) );
  DFFPOSX1 \RF_reg[27][35]  ( .D(n2486), .CLK(clk), .Q(\RF[27][35] ) );
  DFFPOSX1 \RF_reg[27][34]  ( .D(n2485), .CLK(clk), .Q(\RF[27][34] ) );
  DFFPOSX1 \RF_reg[27][33]  ( .D(n2484), .CLK(clk), .Q(\RF[27][33] ) );
  DFFPOSX1 \RF_reg[27][32]  ( .D(n2483), .CLK(clk), .Q(\RF[27][32] ) );
  DFFPOSX1 \RF_reg[27][31]  ( .D(n2482), .CLK(clk), .Q(\RF[27][31] ) );
  DFFPOSX1 \RF_reg[27][30]  ( .D(n2481), .CLK(clk), .Q(\RF[27][30] ) );
  DFFPOSX1 \RF_reg[27][29]  ( .D(n2480), .CLK(clk), .Q(\RF[27][29] ) );
  DFFPOSX1 \RF_reg[27][28]  ( .D(n2479), .CLK(clk), .Q(\RF[27][28] ) );
  DFFPOSX1 \RF_reg[27][27]  ( .D(n2478), .CLK(clk), .Q(\RF[27][27] ) );
  DFFPOSX1 \RF_reg[27][26]  ( .D(n2477), .CLK(clk), .Q(\RF[27][26] ) );
  DFFPOSX1 \RF_reg[27][25]  ( .D(n2476), .CLK(clk), .Q(\RF[27][25] ) );
  DFFPOSX1 \RF_reg[27][24]  ( .D(n2475), .CLK(clk), .Q(\RF[27][24] ) );
  DFFPOSX1 \RF_reg[27][23]  ( .D(n2474), .CLK(clk), .Q(\RF[27][23] ) );
  DFFPOSX1 \RF_reg[27][22]  ( .D(n2473), .CLK(clk), .Q(\RF[27][22] ) );
  DFFPOSX1 \RF_reg[27][21]  ( .D(n2472), .CLK(clk), .Q(\RF[27][21] ) );
  DFFPOSX1 \RF_reg[27][20]  ( .D(n2471), .CLK(clk), .Q(\RF[27][20] ) );
  DFFPOSX1 \RF_reg[27][19]  ( .D(n2470), .CLK(clk), .Q(\RF[27][19] ) );
  DFFPOSX1 \RF_reg[27][18]  ( .D(n2469), .CLK(clk), .Q(\RF[27][18] ) );
  DFFPOSX1 \RF_reg[27][17]  ( .D(n2468), .CLK(clk), .Q(\RF[27][17] ) );
  DFFPOSX1 \RF_reg[27][16]  ( .D(n2467), .CLK(clk), .Q(\RF[27][16] ) );
  DFFPOSX1 \RF_reg[27][15]  ( .D(n2466), .CLK(clk), .Q(\RF[27][15] ) );
  DFFPOSX1 \RF_reg[27][14]  ( .D(n2465), .CLK(clk), .Q(\RF[27][14] ) );
  DFFPOSX1 \RF_reg[27][13]  ( .D(n2464), .CLK(clk), .Q(\RF[27][13] ) );
  DFFPOSX1 \RF_reg[27][12]  ( .D(n2463), .CLK(clk), .Q(\RF[27][12] ) );
  DFFPOSX1 \RF_reg[27][11]  ( .D(n2462), .CLK(clk), .Q(\RF[27][11] ) );
  DFFPOSX1 \RF_reg[27][10]  ( .D(n2461), .CLK(clk), .Q(\RF[27][10] ) );
  DFFPOSX1 \RF_reg[27][9]  ( .D(n2460), .CLK(clk), .Q(\RF[27][9] ) );
  DFFPOSX1 \RF_reg[27][8]  ( .D(n2459), .CLK(clk), .Q(\RF[27][8] ) );
  DFFPOSX1 \RF_reg[27][7]  ( .D(n2458), .CLK(clk), .Q(\RF[27][7] ) );
  DFFPOSX1 \RF_reg[27][6]  ( .D(n2457), .CLK(clk), .Q(\RF[27][6] ) );
  DFFPOSX1 \RF_reg[27][5]  ( .D(n2456), .CLK(clk), .Q(\RF[27][5] ) );
  DFFPOSX1 \RF_reg[27][4]  ( .D(n2455), .CLK(clk), .Q(\RF[27][4] ) );
  DFFPOSX1 \RF_reg[27][3]  ( .D(n2454), .CLK(clk), .Q(\RF[27][3] ) );
  DFFPOSX1 \RF_reg[27][2]  ( .D(n2453), .CLK(clk), .Q(\RF[27][2] ) );
  DFFPOSX1 \RF_reg[27][1]  ( .D(n2452), .CLK(clk), .Q(\RF[27][1] ) );
  DFFPOSX1 \RF_reg[27][0]  ( .D(n2451), .CLK(clk), .Q(\RF[27][0] ) );
  DFFPOSX1 \RF_reg[28][63]  ( .D(n2450), .CLK(clk), .Q(\RF[28][63] ) );
  DFFPOSX1 \RF_reg[28][62]  ( .D(n2449), .CLK(clk), .Q(\RF[28][62] ) );
  DFFPOSX1 \RF_reg[28][61]  ( .D(n2448), .CLK(clk), .Q(\RF[28][61] ) );
  DFFPOSX1 \RF_reg[28][60]  ( .D(n2447), .CLK(clk), .Q(\RF[28][60] ) );
  DFFPOSX1 \RF_reg[28][59]  ( .D(n2446), .CLK(clk), .Q(\RF[28][59] ) );
  DFFPOSX1 \RF_reg[28][58]  ( .D(n2445), .CLK(clk), .Q(\RF[28][58] ) );
  DFFPOSX1 \RF_reg[28][57]  ( .D(n2444), .CLK(clk), .Q(\RF[28][57] ) );
  DFFPOSX1 \RF_reg[28][56]  ( .D(n2443), .CLK(clk), .Q(\RF[28][56] ) );
  DFFPOSX1 \RF_reg[28][55]  ( .D(n2442), .CLK(clk), .Q(\RF[28][55] ) );
  DFFPOSX1 \RF_reg[28][54]  ( .D(n2441), .CLK(clk), .Q(\RF[28][54] ) );
  DFFPOSX1 \RF_reg[28][53]  ( .D(n2440), .CLK(clk), .Q(\RF[28][53] ) );
  DFFPOSX1 \RF_reg[28][52]  ( .D(n2439), .CLK(clk), .Q(\RF[28][52] ) );
  DFFPOSX1 \RF_reg[28][51]  ( .D(n2438), .CLK(clk), .Q(\RF[28][51] ) );
  DFFPOSX1 \RF_reg[28][50]  ( .D(n2437), .CLK(clk), .Q(\RF[28][50] ) );
  DFFPOSX1 \RF_reg[28][49]  ( .D(n2436), .CLK(clk), .Q(\RF[28][49] ) );
  DFFPOSX1 \RF_reg[28][48]  ( .D(n2435), .CLK(clk), .Q(\RF[28][48] ) );
  DFFPOSX1 \RF_reg[28][47]  ( .D(n2434), .CLK(clk), .Q(\RF[28][47] ) );
  DFFPOSX1 \RF_reg[28][46]  ( .D(n2433), .CLK(clk), .Q(\RF[28][46] ) );
  DFFPOSX1 \RF_reg[28][45]  ( .D(n2432), .CLK(clk), .Q(\RF[28][45] ) );
  DFFPOSX1 \RF_reg[28][44]  ( .D(n2431), .CLK(clk), .Q(\RF[28][44] ) );
  DFFPOSX1 \RF_reg[28][43]  ( .D(n2430), .CLK(clk), .Q(\RF[28][43] ) );
  DFFPOSX1 \RF_reg[28][42]  ( .D(n2429), .CLK(clk), .Q(\RF[28][42] ) );
  DFFPOSX1 \RF_reg[28][41]  ( .D(n2428), .CLK(clk), .Q(\RF[28][41] ) );
  DFFPOSX1 \RF_reg[28][40]  ( .D(n2427), .CLK(clk), .Q(\RF[28][40] ) );
  DFFPOSX1 \RF_reg[28][39]  ( .D(n2426), .CLK(clk), .Q(\RF[28][39] ) );
  DFFPOSX1 \RF_reg[28][38]  ( .D(n2425), .CLK(clk), .Q(\RF[28][38] ) );
  DFFPOSX1 \RF_reg[28][37]  ( .D(n2424), .CLK(clk), .Q(\RF[28][37] ) );
  DFFPOSX1 \RF_reg[28][36]  ( .D(n2423), .CLK(clk), .Q(\RF[28][36] ) );
  DFFPOSX1 \RF_reg[28][35]  ( .D(n2422), .CLK(clk), .Q(\RF[28][35] ) );
  DFFPOSX1 \RF_reg[28][34]  ( .D(n2421), .CLK(clk), .Q(\RF[28][34] ) );
  DFFPOSX1 \RF_reg[28][33]  ( .D(n2420), .CLK(clk), .Q(\RF[28][33] ) );
  DFFPOSX1 \RF_reg[28][32]  ( .D(n2419), .CLK(clk), .Q(\RF[28][32] ) );
  DFFPOSX1 \RF_reg[28][31]  ( .D(n2418), .CLK(clk), .Q(\RF[28][31] ) );
  DFFPOSX1 \RF_reg[28][30]  ( .D(n2417), .CLK(clk), .Q(\RF[28][30] ) );
  DFFPOSX1 \RF_reg[28][29]  ( .D(n2416), .CLK(clk), .Q(\RF[28][29] ) );
  DFFPOSX1 \RF_reg[28][28]  ( .D(n2415), .CLK(clk), .Q(\RF[28][28] ) );
  DFFPOSX1 \RF_reg[28][27]  ( .D(n2414), .CLK(clk), .Q(\RF[28][27] ) );
  DFFPOSX1 \RF_reg[28][26]  ( .D(n2413), .CLK(clk), .Q(\RF[28][26] ) );
  DFFPOSX1 \RF_reg[28][25]  ( .D(n2412), .CLK(clk), .Q(\RF[28][25] ) );
  DFFPOSX1 \RF_reg[28][24]  ( .D(n2411), .CLK(clk), .Q(\RF[28][24] ) );
  DFFPOSX1 \RF_reg[28][23]  ( .D(n2410), .CLK(clk), .Q(\RF[28][23] ) );
  DFFPOSX1 \RF_reg[28][22]  ( .D(n2409), .CLK(clk), .Q(\RF[28][22] ) );
  DFFPOSX1 \RF_reg[28][21]  ( .D(n2408), .CLK(clk), .Q(\RF[28][21] ) );
  DFFPOSX1 \RF_reg[28][20]  ( .D(n2407), .CLK(clk), .Q(\RF[28][20] ) );
  DFFPOSX1 \RF_reg[28][19]  ( .D(n2406), .CLK(clk), .Q(\RF[28][19] ) );
  DFFPOSX1 \RF_reg[28][18]  ( .D(n2405), .CLK(clk), .Q(\RF[28][18] ) );
  DFFPOSX1 \RF_reg[28][17]  ( .D(n2404), .CLK(clk), .Q(\RF[28][17] ) );
  DFFPOSX1 \RF_reg[28][16]  ( .D(n2403), .CLK(clk), .Q(\RF[28][16] ) );
  DFFPOSX1 \RF_reg[28][15]  ( .D(n2402), .CLK(clk), .Q(\RF[28][15] ) );
  DFFPOSX1 \RF_reg[28][14]  ( .D(n2401), .CLK(clk), .Q(\RF[28][14] ) );
  DFFPOSX1 \RF_reg[28][13]  ( .D(n2400), .CLK(clk), .Q(\RF[28][13] ) );
  DFFPOSX1 \RF_reg[28][12]  ( .D(n2399), .CLK(clk), .Q(\RF[28][12] ) );
  DFFPOSX1 \RF_reg[28][11]  ( .D(n2398), .CLK(clk), .Q(\RF[28][11] ) );
  DFFPOSX1 \RF_reg[28][10]  ( .D(n2397), .CLK(clk), .Q(\RF[28][10] ) );
  DFFPOSX1 \RF_reg[28][9]  ( .D(n2396), .CLK(clk), .Q(\RF[28][9] ) );
  DFFPOSX1 \RF_reg[28][8]  ( .D(n2395), .CLK(clk), .Q(\RF[28][8] ) );
  DFFPOSX1 \RF_reg[28][7]  ( .D(n2394), .CLK(clk), .Q(\RF[28][7] ) );
  DFFPOSX1 \RF_reg[28][6]  ( .D(n2393), .CLK(clk), .Q(\RF[28][6] ) );
  DFFPOSX1 \RF_reg[28][5]  ( .D(n2392), .CLK(clk), .Q(\RF[28][5] ) );
  DFFPOSX1 \RF_reg[28][4]  ( .D(n2391), .CLK(clk), .Q(\RF[28][4] ) );
  DFFPOSX1 \RF_reg[28][3]  ( .D(n2390), .CLK(clk), .Q(\RF[28][3] ) );
  DFFPOSX1 \RF_reg[28][2]  ( .D(n2389), .CLK(clk), .Q(\RF[28][2] ) );
  DFFPOSX1 \RF_reg[28][1]  ( .D(n2388), .CLK(clk), .Q(\RF[28][1] ) );
  DFFPOSX1 \RF_reg[28][0]  ( .D(n2387), .CLK(clk), .Q(\RF[28][0] ) );
  DFFPOSX1 \RF_reg[29][63]  ( .D(n2386), .CLK(clk), .Q(\RF[29][63] ) );
  DFFPOSX1 \RF_reg[29][62]  ( .D(n2385), .CLK(clk), .Q(\RF[29][62] ) );
  DFFPOSX1 \RF_reg[29][61]  ( .D(n2384), .CLK(clk), .Q(\RF[29][61] ) );
  DFFPOSX1 \RF_reg[29][60]  ( .D(n2383), .CLK(clk), .Q(\RF[29][60] ) );
  DFFPOSX1 \RF_reg[29][59]  ( .D(n2382), .CLK(clk), .Q(\RF[29][59] ) );
  DFFPOSX1 \RF_reg[29][58]  ( .D(n2381), .CLK(clk), .Q(\RF[29][58] ) );
  DFFPOSX1 \RF_reg[29][57]  ( .D(n2380), .CLK(clk), .Q(\RF[29][57] ) );
  DFFPOSX1 \RF_reg[29][56]  ( .D(n2379), .CLK(clk), .Q(\RF[29][56] ) );
  DFFPOSX1 \RF_reg[29][55]  ( .D(n2378), .CLK(clk), .Q(\RF[29][55] ) );
  DFFPOSX1 \RF_reg[29][54]  ( .D(n2377), .CLK(clk), .Q(\RF[29][54] ) );
  DFFPOSX1 \RF_reg[29][53]  ( .D(n2376), .CLK(clk), .Q(\RF[29][53] ) );
  DFFPOSX1 \RF_reg[29][52]  ( .D(n2375), .CLK(clk), .Q(\RF[29][52] ) );
  DFFPOSX1 \RF_reg[29][51]  ( .D(n2374), .CLK(clk), .Q(\RF[29][51] ) );
  DFFPOSX1 \RF_reg[29][50]  ( .D(n2373), .CLK(clk), .Q(\RF[29][50] ) );
  DFFPOSX1 \RF_reg[29][49]  ( .D(n2372), .CLK(clk), .Q(\RF[29][49] ) );
  DFFPOSX1 \RF_reg[29][48]  ( .D(n2371), .CLK(clk), .Q(\RF[29][48] ) );
  DFFPOSX1 \RF_reg[29][47]  ( .D(n2370), .CLK(clk), .Q(\RF[29][47] ) );
  DFFPOSX1 \RF_reg[29][46]  ( .D(n2369), .CLK(clk), .Q(\RF[29][46] ) );
  DFFPOSX1 \RF_reg[29][45]  ( .D(n2368), .CLK(clk), .Q(\RF[29][45] ) );
  DFFPOSX1 \RF_reg[29][44]  ( .D(n2367), .CLK(clk), .Q(\RF[29][44] ) );
  DFFPOSX1 \RF_reg[29][43]  ( .D(n2366), .CLK(clk), .Q(\RF[29][43] ) );
  DFFPOSX1 \RF_reg[29][42]  ( .D(n2365), .CLK(clk), .Q(\RF[29][42] ) );
  DFFPOSX1 \RF_reg[29][41]  ( .D(n2364), .CLK(clk), .Q(\RF[29][41] ) );
  DFFPOSX1 \RF_reg[29][40]  ( .D(n2363), .CLK(clk), .Q(\RF[29][40] ) );
  DFFPOSX1 \RF_reg[29][39]  ( .D(n2362), .CLK(clk), .Q(\RF[29][39] ) );
  DFFPOSX1 \RF_reg[29][38]  ( .D(n2361), .CLK(clk), .Q(\RF[29][38] ) );
  DFFPOSX1 \RF_reg[29][37]  ( .D(n2360), .CLK(clk), .Q(\RF[29][37] ) );
  DFFPOSX1 \RF_reg[29][36]  ( .D(n2359), .CLK(clk), .Q(\RF[29][36] ) );
  DFFPOSX1 \RF_reg[29][35]  ( .D(n2358), .CLK(clk), .Q(\RF[29][35] ) );
  DFFPOSX1 \RF_reg[29][34]  ( .D(n2357), .CLK(clk), .Q(\RF[29][34] ) );
  DFFPOSX1 \RF_reg[29][33]  ( .D(n2356), .CLK(clk), .Q(\RF[29][33] ) );
  DFFPOSX1 \RF_reg[29][32]  ( .D(n2355), .CLK(clk), .Q(\RF[29][32] ) );
  DFFPOSX1 \RF_reg[29][31]  ( .D(n2354), .CLK(clk), .Q(\RF[29][31] ) );
  DFFPOSX1 \RF_reg[29][30]  ( .D(n2353), .CLK(clk), .Q(\RF[29][30] ) );
  DFFPOSX1 \RF_reg[29][29]  ( .D(n2352), .CLK(clk), .Q(\RF[29][29] ) );
  DFFPOSX1 \RF_reg[29][28]  ( .D(n2351), .CLK(clk), .Q(\RF[29][28] ) );
  DFFPOSX1 \RF_reg[29][27]  ( .D(n2350), .CLK(clk), .Q(\RF[29][27] ) );
  DFFPOSX1 \RF_reg[29][26]  ( .D(n2349), .CLK(clk), .Q(\RF[29][26] ) );
  DFFPOSX1 \RF_reg[29][25]  ( .D(n2348), .CLK(clk), .Q(\RF[29][25] ) );
  DFFPOSX1 \RF_reg[29][24]  ( .D(n2347), .CLK(clk), .Q(\RF[29][24] ) );
  DFFPOSX1 \RF_reg[29][23]  ( .D(n2346), .CLK(clk), .Q(\RF[29][23] ) );
  DFFPOSX1 \RF_reg[29][22]  ( .D(n2345), .CLK(clk), .Q(\RF[29][22] ) );
  DFFPOSX1 \RF_reg[29][21]  ( .D(n2344), .CLK(clk), .Q(\RF[29][21] ) );
  DFFPOSX1 \RF_reg[29][20]  ( .D(n2343), .CLK(clk), .Q(\RF[29][20] ) );
  DFFPOSX1 \RF_reg[29][19]  ( .D(n2342), .CLK(clk), .Q(\RF[29][19] ) );
  DFFPOSX1 \RF_reg[29][18]  ( .D(n2341), .CLK(clk), .Q(\RF[29][18] ) );
  DFFPOSX1 \RF_reg[29][17]  ( .D(n2340), .CLK(clk), .Q(\RF[29][17] ) );
  DFFPOSX1 \RF_reg[29][16]  ( .D(n2339), .CLK(clk), .Q(\RF[29][16] ) );
  DFFPOSX1 \RF_reg[29][15]  ( .D(n2338), .CLK(clk), .Q(\RF[29][15] ) );
  DFFPOSX1 \RF_reg[29][14]  ( .D(n2337), .CLK(clk), .Q(\RF[29][14] ) );
  DFFPOSX1 \RF_reg[29][13]  ( .D(n2336), .CLK(clk), .Q(\RF[29][13] ) );
  DFFPOSX1 \RF_reg[29][12]  ( .D(n2335), .CLK(clk), .Q(\RF[29][12] ) );
  DFFPOSX1 \RF_reg[29][11]  ( .D(n2334), .CLK(clk), .Q(\RF[29][11] ) );
  DFFPOSX1 \RF_reg[29][10]  ( .D(n2333), .CLK(clk), .Q(\RF[29][10] ) );
  DFFPOSX1 \RF_reg[29][9]  ( .D(n2332), .CLK(clk), .Q(\RF[29][9] ) );
  DFFPOSX1 \RF_reg[29][8]  ( .D(n2331), .CLK(clk), .Q(\RF[29][8] ) );
  DFFPOSX1 \RF_reg[29][7]  ( .D(n2330), .CLK(clk), .Q(\RF[29][7] ) );
  DFFPOSX1 \RF_reg[29][6]  ( .D(n2329), .CLK(clk), .Q(\RF[29][6] ) );
  DFFPOSX1 \RF_reg[29][5]  ( .D(n2328), .CLK(clk), .Q(\RF[29][5] ) );
  DFFPOSX1 \RF_reg[29][4]  ( .D(n2327), .CLK(clk), .Q(\RF[29][4] ) );
  DFFPOSX1 \RF_reg[29][3]  ( .D(n2326), .CLK(clk), .Q(\RF[29][3] ) );
  DFFPOSX1 \RF_reg[29][2]  ( .D(n2325), .CLK(clk), .Q(\RF[29][2] ) );
  DFFPOSX1 \RF_reg[29][1]  ( .D(n2324), .CLK(clk), .Q(\RF[29][1] ) );
  DFFPOSX1 \RF_reg[29][0]  ( .D(n2323), .CLK(clk), .Q(\RF[29][0] ) );
  DFFPOSX1 \RF_reg[30][63]  ( .D(n2322), .CLK(clk), .Q(\RF[30][63] ) );
  DFFPOSX1 \RF_reg[30][62]  ( .D(n2321), .CLK(clk), .Q(\RF[30][62] ) );
  DFFPOSX1 \RF_reg[30][61]  ( .D(n2320), .CLK(clk), .Q(\RF[30][61] ) );
  DFFPOSX1 \RF_reg[30][60]  ( .D(n2319), .CLK(clk), .Q(\RF[30][60] ) );
  DFFPOSX1 \RF_reg[30][59]  ( .D(n2318), .CLK(clk), .Q(\RF[30][59] ) );
  DFFPOSX1 \RF_reg[30][58]  ( .D(n2317), .CLK(clk), .Q(\RF[30][58] ) );
  DFFPOSX1 \RF_reg[30][57]  ( .D(n2316), .CLK(clk), .Q(\RF[30][57] ) );
  DFFPOSX1 \RF_reg[30][56]  ( .D(n2315), .CLK(clk), .Q(\RF[30][56] ) );
  DFFPOSX1 \RF_reg[30][55]  ( .D(n2314), .CLK(clk), .Q(\RF[30][55] ) );
  DFFPOSX1 \RF_reg[30][54]  ( .D(n2313), .CLK(clk), .Q(\RF[30][54] ) );
  DFFPOSX1 \RF_reg[30][53]  ( .D(n2312), .CLK(clk), .Q(\RF[30][53] ) );
  DFFPOSX1 \RF_reg[30][52]  ( .D(n2311), .CLK(clk), .Q(\RF[30][52] ) );
  DFFPOSX1 \RF_reg[30][51]  ( .D(n2310), .CLK(clk), .Q(\RF[30][51] ) );
  DFFPOSX1 \RF_reg[30][50]  ( .D(n2309), .CLK(clk), .Q(\RF[30][50] ) );
  DFFPOSX1 \RF_reg[30][49]  ( .D(n2308), .CLK(clk), .Q(\RF[30][49] ) );
  DFFPOSX1 \RF_reg[30][48]  ( .D(n2307), .CLK(clk), .Q(\RF[30][48] ) );
  DFFPOSX1 \RF_reg[30][47]  ( .D(n2306), .CLK(clk), .Q(\RF[30][47] ) );
  DFFPOSX1 \RF_reg[30][46]  ( .D(n2305), .CLK(clk), .Q(\RF[30][46] ) );
  DFFPOSX1 \RF_reg[30][45]  ( .D(n2304), .CLK(clk), .Q(\RF[30][45] ) );
  DFFPOSX1 \RF_reg[30][44]  ( .D(n2303), .CLK(clk), .Q(\RF[30][44] ) );
  DFFPOSX1 \RF_reg[30][43]  ( .D(n2302), .CLK(clk), .Q(\RF[30][43] ) );
  DFFPOSX1 \RF_reg[30][42]  ( .D(n2301), .CLK(clk), .Q(\RF[30][42] ) );
  DFFPOSX1 \RF_reg[30][41]  ( .D(n2300), .CLK(clk), .Q(\RF[30][41] ) );
  DFFPOSX1 \RF_reg[30][40]  ( .D(n2299), .CLK(clk), .Q(\RF[30][40] ) );
  DFFPOSX1 \RF_reg[30][39]  ( .D(n2298), .CLK(clk), .Q(\RF[30][39] ) );
  DFFPOSX1 \RF_reg[30][38]  ( .D(n2297), .CLK(clk), .Q(\RF[30][38] ) );
  DFFPOSX1 \RF_reg[30][37]  ( .D(n2296), .CLK(clk), .Q(\RF[30][37] ) );
  DFFPOSX1 \RF_reg[30][36]  ( .D(n2295), .CLK(clk), .Q(\RF[30][36] ) );
  DFFPOSX1 \RF_reg[30][35]  ( .D(n2294), .CLK(clk), .Q(\RF[30][35] ) );
  DFFPOSX1 \RF_reg[30][34]  ( .D(n2293), .CLK(clk), .Q(\RF[30][34] ) );
  DFFPOSX1 \RF_reg[30][33]  ( .D(n2292), .CLK(clk), .Q(\RF[30][33] ) );
  DFFPOSX1 \RF_reg[30][32]  ( .D(n2291), .CLK(clk), .Q(\RF[30][32] ) );
  DFFPOSX1 \RF_reg[30][31]  ( .D(n2290), .CLK(clk), .Q(\RF[30][31] ) );
  DFFPOSX1 \RF_reg[30][30]  ( .D(n2289), .CLK(clk), .Q(\RF[30][30] ) );
  DFFPOSX1 \RF_reg[30][29]  ( .D(n2288), .CLK(clk), .Q(\RF[30][29] ) );
  DFFPOSX1 \RF_reg[30][28]  ( .D(n2287), .CLK(clk), .Q(\RF[30][28] ) );
  DFFPOSX1 \RF_reg[30][27]  ( .D(n2286), .CLK(clk), .Q(\RF[30][27] ) );
  DFFPOSX1 \RF_reg[30][26]  ( .D(n2285), .CLK(clk), .Q(\RF[30][26] ) );
  DFFPOSX1 \RF_reg[30][25]  ( .D(n2284), .CLK(clk), .Q(\RF[30][25] ) );
  DFFPOSX1 \RF_reg[30][24]  ( .D(n2283), .CLK(clk), .Q(\RF[30][24] ) );
  DFFPOSX1 \RF_reg[30][23]  ( .D(n2282), .CLK(clk), .Q(\RF[30][23] ) );
  DFFPOSX1 \RF_reg[30][22]  ( .D(n2281), .CLK(clk), .Q(\RF[30][22] ) );
  DFFPOSX1 \RF_reg[30][21]  ( .D(n2280), .CLK(clk), .Q(\RF[30][21] ) );
  DFFPOSX1 \RF_reg[30][20]  ( .D(n2279), .CLK(clk), .Q(\RF[30][20] ) );
  DFFPOSX1 \RF_reg[30][19]  ( .D(n2278), .CLK(clk), .Q(\RF[30][19] ) );
  DFFPOSX1 \RF_reg[30][18]  ( .D(n2277), .CLK(clk), .Q(\RF[30][18] ) );
  DFFPOSX1 \RF_reg[30][17]  ( .D(n2276), .CLK(clk), .Q(\RF[30][17] ) );
  DFFPOSX1 \RF_reg[30][16]  ( .D(n2275), .CLK(clk), .Q(\RF[30][16] ) );
  DFFPOSX1 \RF_reg[30][15]  ( .D(n2274), .CLK(clk), .Q(\RF[30][15] ) );
  DFFPOSX1 \RF_reg[30][14]  ( .D(n2273), .CLK(clk), .Q(\RF[30][14] ) );
  DFFPOSX1 \RF_reg[30][13]  ( .D(n2272), .CLK(clk), .Q(\RF[30][13] ) );
  DFFPOSX1 \RF_reg[30][12]  ( .D(n2271), .CLK(clk), .Q(\RF[30][12] ) );
  DFFPOSX1 \RF_reg[30][11]  ( .D(n2270), .CLK(clk), .Q(\RF[30][11] ) );
  DFFPOSX1 \RF_reg[30][10]  ( .D(n2269), .CLK(clk), .Q(\RF[30][10] ) );
  DFFPOSX1 \RF_reg[30][9]  ( .D(n2268), .CLK(clk), .Q(\RF[30][9] ) );
  DFFPOSX1 \RF_reg[30][8]  ( .D(n2267), .CLK(clk), .Q(\RF[30][8] ) );
  DFFPOSX1 \RF_reg[30][7]  ( .D(n2266), .CLK(clk), .Q(\RF[30][7] ) );
  DFFPOSX1 \RF_reg[30][6]  ( .D(n2265), .CLK(clk), .Q(\RF[30][6] ) );
  DFFPOSX1 \RF_reg[30][5]  ( .D(n2264), .CLK(clk), .Q(\RF[30][5] ) );
  DFFPOSX1 \RF_reg[30][4]  ( .D(n2263), .CLK(clk), .Q(\RF[30][4] ) );
  DFFPOSX1 \RF_reg[30][3]  ( .D(n2262), .CLK(clk), .Q(\RF[30][3] ) );
  DFFPOSX1 \RF_reg[30][2]  ( .D(n2261), .CLK(clk), .Q(\RF[30][2] ) );
  DFFPOSX1 \RF_reg[30][1]  ( .D(n2260), .CLK(clk), .Q(\RF[30][1] ) );
  DFFPOSX1 \RF_reg[30][0]  ( .D(n2259), .CLK(clk), .Q(\RF[30][0] ) );
  DFFPOSX1 \RF_reg[31][63]  ( .D(n2258), .CLK(clk), .Q(\RF[31][63] ) );
  DFFPOSX1 \RF_reg[31][62]  ( .D(n2257), .CLK(clk), .Q(\RF[31][62] ) );
  DFFPOSX1 \RF_reg[31][61]  ( .D(n2256), .CLK(clk), .Q(\RF[31][61] ) );
  DFFPOSX1 \RF_reg[31][60]  ( .D(n2255), .CLK(clk), .Q(\RF[31][60] ) );
  DFFPOSX1 \RF_reg[31][59]  ( .D(n2254), .CLK(clk), .Q(\RF[31][59] ) );
  DFFPOSX1 \RF_reg[31][58]  ( .D(n2253), .CLK(clk), .Q(\RF[31][58] ) );
  DFFPOSX1 \RF_reg[31][57]  ( .D(n2252), .CLK(clk), .Q(\RF[31][57] ) );
  DFFPOSX1 \RF_reg[31][56]  ( .D(n2251), .CLK(clk), .Q(\RF[31][56] ) );
  DFFPOSX1 \RF_reg[31][55]  ( .D(n2250), .CLK(clk), .Q(\RF[31][55] ) );
  DFFPOSX1 \RF_reg[31][54]  ( .D(n2249), .CLK(clk), .Q(\RF[31][54] ) );
  DFFPOSX1 \RF_reg[31][53]  ( .D(n2248), .CLK(clk), .Q(\RF[31][53] ) );
  DFFPOSX1 \RF_reg[31][52]  ( .D(n2247), .CLK(clk), .Q(\RF[31][52] ) );
  DFFPOSX1 \RF_reg[31][51]  ( .D(n2246), .CLK(clk), .Q(\RF[31][51] ) );
  DFFPOSX1 \RF_reg[31][50]  ( .D(n2245), .CLK(clk), .Q(\RF[31][50] ) );
  DFFPOSX1 \RF_reg[31][49]  ( .D(n2244), .CLK(clk), .Q(\RF[31][49] ) );
  DFFPOSX1 \RF_reg[31][48]  ( .D(n2243), .CLK(clk), .Q(\RF[31][48] ) );
  DFFPOSX1 \RF_reg[31][47]  ( .D(n2242), .CLK(clk), .Q(\RF[31][47] ) );
  DFFPOSX1 \RF_reg[31][46]  ( .D(n2241), .CLK(clk), .Q(\RF[31][46] ) );
  DFFPOSX1 \RF_reg[31][45]  ( .D(n2240), .CLK(clk), .Q(\RF[31][45] ) );
  DFFPOSX1 \RF_reg[31][44]  ( .D(n2239), .CLK(clk), .Q(\RF[31][44] ) );
  DFFPOSX1 \RF_reg[31][43]  ( .D(n2238), .CLK(clk), .Q(\RF[31][43] ) );
  DFFPOSX1 \RF_reg[31][42]  ( .D(n2237), .CLK(clk), .Q(\RF[31][42] ) );
  DFFPOSX1 \RF_reg[31][41]  ( .D(n2236), .CLK(clk), .Q(\RF[31][41] ) );
  DFFPOSX1 \RF_reg[31][40]  ( .D(n2235), .CLK(clk), .Q(\RF[31][40] ) );
  DFFPOSX1 \RF_reg[31][39]  ( .D(n2234), .CLK(clk), .Q(\RF[31][39] ) );
  DFFPOSX1 \RF_reg[31][38]  ( .D(n2233), .CLK(clk), .Q(\RF[31][38] ) );
  DFFPOSX1 \RF_reg[31][37]  ( .D(n2232), .CLK(clk), .Q(\RF[31][37] ) );
  DFFPOSX1 \RF_reg[31][36]  ( .D(n2231), .CLK(clk), .Q(\RF[31][36] ) );
  DFFPOSX1 \RF_reg[31][35]  ( .D(n2230), .CLK(clk), .Q(\RF[31][35] ) );
  DFFPOSX1 \RF_reg[31][34]  ( .D(n2229), .CLK(clk), .Q(\RF[31][34] ) );
  DFFPOSX1 \RF_reg[31][33]  ( .D(n2228), .CLK(clk), .Q(\RF[31][33] ) );
  DFFPOSX1 \RF_reg[31][32]  ( .D(n2227), .CLK(clk), .Q(\RF[31][32] ) );
  DFFPOSX1 \RF_reg[31][31]  ( .D(n2226), .CLK(clk), .Q(\RF[31][31] ) );
  DFFPOSX1 \RF_reg[31][30]  ( .D(n2225), .CLK(clk), .Q(\RF[31][30] ) );
  DFFPOSX1 \RF_reg[31][29]  ( .D(n2224), .CLK(clk), .Q(\RF[31][29] ) );
  DFFPOSX1 \RF_reg[31][28]  ( .D(n2223), .CLK(clk), .Q(\RF[31][28] ) );
  DFFPOSX1 \RF_reg[31][27]  ( .D(n2222), .CLK(clk), .Q(\RF[31][27] ) );
  DFFPOSX1 \RF_reg[31][26]  ( .D(n2221), .CLK(clk), .Q(\RF[31][26] ) );
  DFFPOSX1 \RF_reg[31][25]  ( .D(n2220), .CLK(clk), .Q(\RF[31][25] ) );
  DFFPOSX1 \RF_reg[31][24]  ( .D(n2219), .CLK(clk), .Q(\RF[31][24] ) );
  DFFPOSX1 \RF_reg[31][23]  ( .D(n2218), .CLK(clk), .Q(\RF[31][23] ) );
  DFFPOSX1 \RF_reg[31][22]  ( .D(n2217), .CLK(clk), .Q(\RF[31][22] ) );
  DFFPOSX1 \RF_reg[31][21]  ( .D(n2216), .CLK(clk), .Q(\RF[31][21] ) );
  DFFPOSX1 \RF_reg[31][20]  ( .D(n2215), .CLK(clk), .Q(\RF[31][20] ) );
  DFFPOSX1 \RF_reg[31][19]  ( .D(n2214), .CLK(clk), .Q(\RF[31][19] ) );
  DFFPOSX1 \RF_reg[31][18]  ( .D(n2213), .CLK(clk), .Q(\RF[31][18] ) );
  DFFPOSX1 \RF_reg[31][17]  ( .D(n2212), .CLK(clk), .Q(\RF[31][17] ) );
  DFFPOSX1 \RF_reg[31][16]  ( .D(n2211), .CLK(clk), .Q(\RF[31][16] ) );
  DFFPOSX1 \RF_reg[31][15]  ( .D(n2210), .CLK(clk), .Q(\RF[31][15] ) );
  DFFPOSX1 \RF_reg[31][14]  ( .D(n2209), .CLK(clk), .Q(\RF[31][14] ) );
  DFFPOSX1 \RF_reg[31][13]  ( .D(n2208), .CLK(clk), .Q(\RF[31][13] ) );
  DFFPOSX1 \RF_reg[31][12]  ( .D(n2207), .CLK(clk), .Q(\RF[31][12] ) );
  DFFPOSX1 \RF_reg[31][11]  ( .D(n2206), .CLK(clk), .Q(\RF[31][11] ) );
  DFFPOSX1 \RF_reg[31][10]  ( .D(n2205), .CLK(clk), .Q(\RF[31][10] ) );
  DFFPOSX1 \RF_reg[31][9]  ( .D(n2204), .CLK(clk), .Q(\RF[31][9] ) );
  DFFPOSX1 \RF_reg[31][8]  ( .D(n2203), .CLK(clk), .Q(\RF[31][8] ) );
  DFFPOSX1 \RF_reg[31][7]  ( .D(n2202), .CLK(clk), .Q(\RF[31][7] ) );
  DFFPOSX1 \RF_reg[31][6]  ( .D(n2201), .CLK(clk), .Q(\RF[31][6] ) );
  DFFPOSX1 \RF_reg[31][5]  ( .D(n2200), .CLK(clk), .Q(\RF[31][5] ) );
  DFFPOSX1 \RF_reg[31][4]  ( .D(n2199), .CLK(clk), .Q(\RF[31][4] ) );
  DFFPOSX1 \RF_reg[31][3]  ( .D(n2198), .CLK(clk), .Q(\RF[31][3] ) );
  DFFPOSX1 \RF_reg[31][2]  ( .D(n2197), .CLK(clk), .Q(\RF[31][2] ) );
  DFFPOSX1 \RF_reg[31][1]  ( .D(n2196), .CLK(clk), .Q(\RF[31][1] ) );
  DFFPOSX1 \RF_reg[31][0]  ( .D(n2195), .CLK(clk), .Q(\RF[31][0] ) );
  OAI21X1 U169 ( .A(n10763), .B(n10830), .C(n6301), .Y(n2195) );
  OAI21X1 U171 ( .A(n10763), .B(n10829), .C(n6300), .Y(n2196) );
  OAI21X1 U173 ( .A(n10763), .B(n10828), .C(n6169), .Y(n2197) );
  OAI21X1 U175 ( .A(n10763), .B(n10827), .C(n6037), .Y(n2198) );
  OAI21X1 U177 ( .A(n10763), .B(n10826), .C(n5905), .Y(n2199) );
  OAI21X1 U179 ( .A(n10763), .B(n10825), .C(n5770), .Y(n2200) );
  OAI21X1 U181 ( .A(n10763), .B(n10824), .C(n5652), .Y(n2201) );
  OAI21X1 U183 ( .A(n10763), .B(n10823), .C(n5534), .Y(n2202) );
  OAI21X1 U185 ( .A(n10763), .B(n10822), .C(n5416), .Y(n2203) );
  OAI21X1 U187 ( .A(n10763), .B(n10821), .C(n5298), .Y(n2204) );
  OAI21X1 U189 ( .A(n10763), .B(n10820), .C(n5189), .Y(n2205) );
  OAI21X1 U191 ( .A(n10763), .B(n10819), .C(n5080), .Y(n2206) );
  OAI21X1 U193 ( .A(n10763), .B(n10818), .C(n4971), .Y(n2207) );
  OAI21X1 U195 ( .A(n10763), .B(n10817), .C(n6299), .Y(n2208) );
  OAI21X1 U197 ( .A(n10763), .B(n10816), .C(n6168), .Y(n2209) );
  OAI21X1 U199 ( .A(n10763), .B(n10815), .C(n6036), .Y(n2210) );
  OAI21X1 U201 ( .A(n10764), .B(n10814), .C(n5904), .Y(n2211) );
  OAI21X1 U203 ( .A(n10764), .B(n10813), .C(n5769), .Y(n2212) );
  OAI21X1 U205 ( .A(n10763), .B(n10812), .C(n5651), .Y(n2213) );
  OAI21X1 U207 ( .A(n10764), .B(n10811), .C(n5533), .Y(n2214) );
  OAI21X1 U209 ( .A(n10764), .B(n10810), .C(n5415), .Y(n2215) );
  OAI21X1 U211 ( .A(n10764), .B(n10809), .C(n5297), .Y(n2216) );
  OAI21X1 U213 ( .A(n10764), .B(n10808), .C(n5188), .Y(n2217) );
  OAI21X1 U215 ( .A(n10763), .B(n10807), .C(n5079), .Y(n2218) );
  OAI21X1 U217 ( .A(n10763), .B(n10806), .C(n4862), .Y(n2219) );
  OAI21X1 U219 ( .A(n10763), .B(n10805), .C(n5414), .Y(n2220) );
  OAI21X1 U221 ( .A(n10763), .B(n10804), .C(n6167), .Y(n2221) );
  OAI21X1 U223 ( .A(n10763), .B(n10803), .C(n6035), .Y(n2222) );
  OAI21X1 U225 ( .A(n10764), .B(n10802), .C(n5903), .Y(n2223) );
  OAI21X1 U227 ( .A(n10763), .B(n10801), .C(n5768), .Y(n2224) );
  OAI21X1 U229 ( .A(n10764), .B(n10800), .C(n5650), .Y(n2225) );
  OAI21X1 U231 ( .A(n10763), .B(n10799), .C(n5532), .Y(n2226) );
  OAI21X1 U233 ( .A(n10763), .B(n10798), .C(n6298), .Y(n2227) );
  OAI21X1 U235 ( .A(n10763), .B(n10797), .C(n5296), .Y(n2228) );
  OAI21X1 U237 ( .A(n10764), .B(n10796), .C(n5187), .Y(n2229) );
  OAI21X1 U239 ( .A(n10763), .B(n10795), .C(n5078), .Y(n2230) );
  OAI21X1 U241 ( .A(n10763), .B(n10794), .C(n4970), .Y(n2231) );
  OAI21X1 U243 ( .A(n10764), .B(n10793), .C(n6166), .Y(n2232) );
  OAI21X1 U245 ( .A(n10763), .B(n10792), .C(n5649), .Y(n2233) );
  OAI21X1 U247 ( .A(n10763), .B(n10791), .C(n6034), .Y(n2234) );
  OAI21X1 U249 ( .A(n10763), .B(n10790), .C(n5902), .Y(n2235) );
  OAI21X1 U251 ( .A(n10764), .B(n10789), .C(n5767), .Y(n2236) );
  OAI21X1 U253 ( .A(n10764), .B(n10788), .C(n4969), .Y(n2237) );
  OAI21X1 U255 ( .A(n10763), .B(n10787), .C(n5531), .Y(n2238) );
  OAI21X1 U257 ( .A(n10764), .B(n10786), .C(n5295), .Y(n2239) );
  OAI21X1 U259 ( .A(n10764), .B(n10785), .C(n6297), .Y(n2240) );
  OAI21X1 U261 ( .A(n10763), .B(n10784), .C(n4861), .Y(n2241) );
  OAI21X1 U263 ( .A(n10763), .B(n10783), .C(n5413), .Y(n2242) );
  OAI21X1 U265 ( .A(n10763), .B(n10782), .C(n4755), .Y(n2243) );
  OAI21X1 U267 ( .A(n10764), .B(n10781), .C(n4648), .Y(n2244) );
  OAI21X1 U269 ( .A(n10764), .B(n10780), .C(n4541), .Y(n2245) );
  OAI21X1 U271 ( .A(n10763), .B(n10779), .C(n4434), .Y(n2246) );
  OAI21X1 U273 ( .A(n10764), .B(n10778), .C(n4433), .Y(n2247) );
  OAI21X1 U275 ( .A(n10764), .B(n10777), .C(n4647), .Y(n2248) );
  OAI21X1 U277 ( .A(n10763), .B(n10776), .C(n4432), .Y(n2249) );
  OAI21X1 U279 ( .A(n10764), .B(n10775), .C(n4431), .Y(n2250) );
  OAI21X1 U281 ( .A(n10764), .B(n10774), .C(n5077), .Y(n2251) );
  OAI21X1 U283 ( .A(n10763), .B(n10773), .C(n4860), .Y(n2252) );
  OAI21X1 U285 ( .A(n10764), .B(n10772), .C(n4754), .Y(n2253) );
  OAI21X1 U287 ( .A(n10763), .B(n10771), .C(n4968), .Y(n2254) );
  OAI21X1 U289 ( .A(n10763), .B(n10770), .C(n4430), .Y(n2255) );
  OAI21X1 U291 ( .A(n10763), .B(n10769), .C(n4646), .Y(n2256) );
  OAI21X1 U293 ( .A(n10764), .B(n10768), .C(n4429), .Y(n2257) );
  OAI21X1 U295 ( .A(n10764), .B(n10767), .C(n5186), .Y(n2258) );
  OAI21X1 U297 ( .A(n5906), .B(n5774), .C(reset_n), .Y(n166) );
  OAI21X1 U298 ( .A(n10761), .B(n10830), .C(n6165), .Y(n2259) );
  OAI21X1 U300 ( .A(n10761), .B(n10829), .C(n6164), .Y(n2260) );
  OAI21X1 U302 ( .A(n10761), .B(n10828), .C(n6296), .Y(n2261) );
  OAI21X1 U304 ( .A(n10761), .B(n10827), .C(n5901), .Y(n2262) );
  OAI21X1 U306 ( .A(n10761), .B(n10826), .C(n6033), .Y(n2263) );
  OAI21X1 U308 ( .A(n10761), .B(n10825), .C(n5648), .Y(n2264) );
  OAI21X1 U310 ( .A(n10761), .B(n10824), .C(n5766), .Y(n2265) );
  OAI21X1 U312 ( .A(n10761), .B(n10823), .C(n5412), .Y(n2266) );
  OAI21X1 U314 ( .A(n10761), .B(n10822), .C(n5530), .Y(n2267) );
  OAI21X1 U316 ( .A(n10761), .B(n10821), .C(n5185), .Y(n2268) );
  OAI21X1 U318 ( .A(n10761), .B(n10820), .C(n5294), .Y(n2269) );
  OAI21X1 U320 ( .A(n10761), .B(n10819), .C(n4967), .Y(n2270) );
  OAI21X1 U322 ( .A(n10761), .B(n10818), .C(n5076), .Y(n2271) );
  OAI21X1 U324 ( .A(n10761), .B(n10817), .C(n6163), .Y(n2272) );
  OAI21X1 U326 ( .A(n10761), .B(n10816), .C(n6295), .Y(n2273) );
  OAI21X1 U328 ( .A(n10761), .B(n10815), .C(n5900), .Y(n2274) );
  OAI21X1 U330 ( .A(n10762), .B(n10814), .C(n6032), .Y(n2275) );
  OAI21X1 U332 ( .A(n10762), .B(n10813), .C(n5647), .Y(n2276) );
  OAI21X1 U334 ( .A(n10761), .B(n10812), .C(n5765), .Y(n2277) );
  OAI21X1 U336 ( .A(n10762), .B(n10811), .C(n5411), .Y(n2278) );
  OAI21X1 U338 ( .A(n10762), .B(n10810), .C(n5529), .Y(n2279) );
  OAI21X1 U340 ( .A(n10762), .B(n10809), .C(n5184), .Y(n2280) );
  OAI21X1 U342 ( .A(n10762), .B(n10808), .C(n5293), .Y(n2281) );
  OAI21X1 U344 ( .A(n10761), .B(n10807), .C(n4966), .Y(n2282) );
  OAI21X1 U346 ( .A(n10761), .B(n10806), .C(n4753), .Y(n2283) );
  OAI21X1 U348 ( .A(n10761), .B(n10805), .C(n5528), .Y(n2284) );
  OAI21X1 U350 ( .A(n10761), .B(n10804), .C(n6294), .Y(n2285) );
  OAI21X1 U352 ( .A(n10761), .B(n10803), .C(n5899), .Y(n2286) );
  OAI21X1 U354 ( .A(n10762), .B(n10802), .C(n6031), .Y(n2287) );
  OAI21X1 U356 ( .A(n10761), .B(n10801), .C(n5646), .Y(n2288) );
  OAI21X1 U358 ( .A(n10762), .B(n10800), .C(n5764), .Y(n2289) );
  OAI21X1 U360 ( .A(n10761), .B(n10799), .C(n5410), .Y(n2290) );
  OAI21X1 U362 ( .A(n10761), .B(n10798), .C(n6162), .Y(n2291) );
  OAI21X1 U364 ( .A(n10761), .B(n10797), .C(n5183), .Y(n2292) );
  OAI21X1 U366 ( .A(n10762), .B(n10796), .C(n5292), .Y(n2293) );
  OAI21X1 U368 ( .A(n10761), .B(n10795), .C(n4965), .Y(n2294) );
  OAI21X1 U370 ( .A(n10761), .B(n10794), .C(n5075), .Y(n2295) );
  OAI21X1 U372 ( .A(n10762), .B(n10793), .C(n6293), .Y(n2296) );
  OAI21X1 U374 ( .A(n10761), .B(n10792), .C(n5763), .Y(n2297) );
  OAI21X1 U376 ( .A(n10761), .B(n10791), .C(n5898), .Y(n2298) );
  OAI21X1 U378 ( .A(n10761), .B(n10790), .C(n6030), .Y(n2299) );
  OAI21X1 U380 ( .A(n10762), .B(n10789), .C(n5645), .Y(n2300) );
  OAI21X1 U382 ( .A(n10762), .B(n10788), .C(n5074), .Y(n2301) );
  OAI21X1 U384 ( .A(n10761), .B(n10787), .C(n5409), .Y(n2302) );
  OAI21X1 U386 ( .A(n10762), .B(n10786), .C(n5182), .Y(n2303) );
  OAI21X1 U388 ( .A(n10762), .B(n10785), .C(n6161), .Y(n2304) );
  OAI21X1 U390 ( .A(n10761), .B(n10784), .C(n4752), .Y(n2305) );
  OAI21X1 U392 ( .A(n10761), .B(n10783), .C(n5527), .Y(n2306) );
  OAI21X1 U394 ( .A(n10761), .B(n10782), .C(n4859), .Y(n2307) );
  OAI21X1 U396 ( .A(n10762), .B(n10781), .C(n4540), .Y(n2308) );
  OAI21X1 U398 ( .A(n10762), .B(n10780), .C(n4645), .Y(n2309) );
  OAI21X1 U400 ( .A(n10761), .B(n10779), .C(n4428), .Y(n2310) );
  OAI21X1 U402 ( .A(n10762), .B(n10778), .C(n4427), .Y(n2311) );
  OAI21X1 U404 ( .A(n10762), .B(n10777), .C(n4539), .Y(n2312) );
  OAI21X1 U406 ( .A(n10761), .B(n10776), .C(n4426), .Y(n2313) );
  OAI21X1 U408 ( .A(n10762), .B(n10775), .C(n4425), .Y(n2314) );
  OAI21X1 U410 ( .A(n10762), .B(n10774), .C(n4964), .Y(n2315) );
  OAI21X1 U412 ( .A(n10761), .B(n10773), .C(n4751), .Y(n2316) );
  OAI21X1 U414 ( .A(n10762), .B(n10772), .C(n4858), .Y(n2317) );
  OAI21X1 U416 ( .A(n10761), .B(n10771), .C(n5073), .Y(n2318) );
  OAI21X1 U418 ( .A(n10761), .B(n10770), .C(n4424), .Y(n2319) );
  OAI21X1 U420 ( .A(n10761), .B(n10769), .C(n4538), .Y(n2320) );
  OAI21X1 U422 ( .A(n10762), .B(n10768), .C(n4423), .Y(n2321) );
  OAI21X1 U424 ( .A(n10762), .B(n10767), .C(n5291), .Y(n2322) );
  OAI21X1 U426 ( .A(n5906), .B(n5773), .C(reset_n), .Y(n233) );
  OAI21X1 U427 ( .A(n10759), .B(n10830), .C(n6029), .Y(n2323) );
  OAI21X1 U429 ( .A(n10759), .B(n10829), .C(n6028), .Y(n2324) );
  OAI21X1 U431 ( .A(n10759), .B(n10828), .C(n5897), .Y(n2325) );
  OAI21X1 U433 ( .A(n10759), .B(n10827), .C(n6292), .Y(n2326) );
  OAI21X1 U435 ( .A(n10759), .B(n10826), .C(n6160), .Y(n2327) );
  OAI21X1 U437 ( .A(n10759), .B(n10825), .C(n5526), .Y(n2328) );
  OAI21X1 U439 ( .A(n10759), .B(n10824), .C(n5408), .Y(n2329) );
  OAI21X1 U441 ( .A(n10759), .B(n10823), .C(n5762), .Y(n2330) );
  OAI21X1 U443 ( .A(n10759), .B(n10822), .C(n5644), .Y(n2331) );
  OAI21X1 U445 ( .A(n10759), .B(n10821), .C(n5072), .Y(n2332) );
  OAI21X1 U447 ( .A(n10759), .B(n10820), .C(n4963), .Y(n2333) );
  OAI21X1 U449 ( .A(n10759), .B(n10819), .C(n5290), .Y(n2334) );
  OAI21X1 U451 ( .A(n10759), .B(n10818), .C(n5181), .Y(n2335) );
  OAI21X1 U453 ( .A(n10759), .B(n10817), .C(n6027), .Y(n2336) );
  OAI21X1 U455 ( .A(n10759), .B(n10816), .C(n5896), .Y(n2337) );
  OAI21X1 U457 ( .A(n10759), .B(n10815), .C(n6291), .Y(n2338) );
  OAI21X1 U459 ( .A(n10760), .B(n10814), .C(n6159), .Y(n2339) );
  OAI21X1 U461 ( .A(n10760), .B(n10813), .C(n5525), .Y(n2340) );
  OAI21X1 U463 ( .A(n10759), .B(n10812), .C(n5407), .Y(n2341) );
  OAI21X1 U465 ( .A(n10760), .B(n10811), .C(n5761), .Y(n2342) );
  OAI21X1 U467 ( .A(n10760), .B(n10810), .C(n5643), .Y(n2343) );
  OAI21X1 U469 ( .A(n10760), .B(n10809), .C(n5071), .Y(n2344) );
  OAI21X1 U471 ( .A(n10760), .B(n10808), .C(n4962), .Y(n2345) );
  OAI21X1 U473 ( .A(n10759), .B(n10807), .C(n5289), .Y(n2346) );
  OAI21X1 U475 ( .A(n10759), .B(n10806), .C(n4644), .Y(n2347) );
  OAI21X1 U477 ( .A(n10759), .B(n10805), .C(n5642), .Y(n2348) );
  OAI21X1 U479 ( .A(n10759), .B(n10804), .C(n5895), .Y(n2349) );
  OAI21X1 U481 ( .A(n10759), .B(n10803), .C(n6290), .Y(n2350) );
  OAI21X1 U483 ( .A(n10760), .B(n10802), .C(n6158), .Y(n2351) );
  OAI21X1 U485 ( .A(n10759), .B(n10801), .C(n5524), .Y(n2352) );
  OAI21X1 U487 ( .A(n10760), .B(n10800), .C(n5406), .Y(n2353) );
  OAI21X1 U489 ( .A(n10759), .B(n10799), .C(n5760), .Y(n2354) );
  OAI21X1 U491 ( .A(n10759), .B(n10798), .C(n6026), .Y(n2355) );
  OAI21X1 U493 ( .A(n10759), .B(n10797), .C(n5070), .Y(n2356) );
  OAI21X1 U495 ( .A(n10760), .B(n10796), .C(n4961), .Y(n2357) );
  OAI21X1 U497 ( .A(n10759), .B(n10795), .C(n5288), .Y(n2358) );
  OAI21X1 U499 ( .A(n10759), .B(n10794), .C(n5180), .Y(n2359) );
  OAI21X1 U501 ( .A(n10760), .B(n10793), .C(n5894), .Y(n2360) );
  OAI21X1 U503 ( .A(n10759), .B(n10792), .C(n5405), .Y(n2361) );
  OAI21X1 U505 ( .A(n10759), .B(n10791), .C(n6289), .Y(n2362) );
  OAI21X1 U507 ( .A(n10759), .B(n10790), .C(n6157), .Y(n2363) );
  OAI21X1 U509 ( .A(n10760), .B(n10789), .C(n5523), .Y(n2364) );
  OAI21X1 U511 ( .A(n10760), .B(n10788), .C(n5179), .Y(n2365) );
  OAI21X1 U513 ( .A(n10759), .B(n10787), .C(n5759), .Y(n2366) );
  OAI21X1 U515 ( .A(n10760), .B(n10786), .C(n5069), .Y(n2367) );
  OAI21X1 U517 ( .A(n10760), .B(n10785), .C(n6025), .Y(n2368) );
  OAI21X1 U519 ( .A(n10759), .B(n10784), .C(n4643), .Y(n2369) );
  OAI21X1 U521 ( .A(n10759), .B(n10783), .C(n5641), .Y(n2370) );
  OAI21X1 U523 ( .A(n10759), .B(n10782), .C(n4537), .Y(n2371) );
  OAI21X1 U525 ( .A(n10760), .B(n10781), .C(n4857), .Y(n2372) );
  OAI21X1 U527 ( .A(n10760), .B(n10780), .C(n4750), .Y(n2373) );
  OAI21X1 U529 ( .A(n10759), .B(n10779), .C(n4422), .Y(n2374) );
  OAI21X1 U531 ( .A(n10760), .B(n10778), .C(n4421), .Y(n2375) );
  OAI21X1 U533 ( .A(n10760), .B(n10777), .C(n4856), .Y(n2376) );
  OAI21X1 U535 ( .A(n10759), .B(n10776), .C(n4420), .Y(n2377) );
  OAI21X1 U537 ( .A(n10760), .B(n10775), .C(n4419), .Y(n2378) );
  OAI21X1 U539 ( .A(n10760), .B(n10774), .C(n5287), .Y(n2379) );
  OAI21X1 U541 ( .A(n10759), .B(n10773), .C(n4642), .Y(n2380) );
  OAI21X1 U543 ( .A(n10760), .B(n10772), .C(n4536), .Y(n2381) );
  OAI21X1 U545 ( .A(n10759), .B(n10771), .C(n5178), .Y(n2382) );
  OAI21X1 U547 ( .A(n10759), .B(n10770), .C(n4418), .Y(n2383) );
  OAI21X1 U549 ( .A(n10759), .B(n10769), .C(n4855), .Y(n2384) );
  OAI21X1 U551 ( .A(n10760), .B(n10768), .C(n4417), .Y(n2385) );
  OAI21X1 U553 ( .A(n10760), .B(n10767), .C(n4960), .Y(n2386) );
  OAI21X1 U555 ( .A(n5906), .B(n5772), .C(reset_n), .Y(n299) );
  OAI21X1 U556 ( .A(n10757), .B(n10830), .C(n5893), .Y(n2387) );
  OAI21X1 U558 ( .A(n10757), .B(n10829), .C(n5892), .Y(n2388) );
  OAI21X1 U560 ( .A(n10757), .B(n10828), .C(n6024), .Y(n2389) );
  OAI21X1 U562 ( .A(n10757), .B(n10827), .C(n6156), .Y(n2390) );
  OAI21X1 U564 ( .A(n10757), .B(n10826), .C(n6288), .Y(n2391) );
  OAI21X1 U566 ( .A(n10757), .B(n10825), .C(n5404), .Y(n2392) );
  OAI21X1 U568 ( .A(n10757), .B(n10824), .C(n5522), .Y(n2393) );
  OAI21X1 U570 ( .A(n10757), .B(n10823), .C(n5640), .Y(n2394) );
  OAI21X1 U572 ( .A(n10757), .B(n10822), .C(n5758), .Y(n2395) );
  OAI21X1 U574 ( .A(n10757), .B(n10821), .C(n4959), .Y(n2396) );
  OAI21X1 U576 ( .A(n10757), .B(n10820), .C(n5068), .Y(n2397) );
  OAI21X1 U578 ( .A(n10757), .B(n10819), .C(n5177), .Y(n2398) );
  OAI21X1 U580 ( .A(n10757), .B(n10818), .C(n5286), .Y(n2399) );
  OAI21X1 U582 ( .A(n10757), .B(n10817), .C(n5891), .Y(n2400) );
  OAI21X1 U584 ( .A(n10757), .B(n10816), .C(n6023), .Y(n2401) );
  OAI21X1 U586 ( .A(n10757), .B(n10815), .C(n6155), .Y(n2402) );
  OAI21X1 U588 ( .A(n10758), .B(n10814), .C(n6287), .Y(n2403) );
  OAI21X1 U590 ( .A(n10758), .B(n10813), .C(n5403), .Y(n2404) );
  OAI21X1 U592 ( .A(n10757), .B(n10812), .C(n5521), .Y(n2405) );
  OAI21X1 U594 ( .A(n10758), .B(n10811), .C(n5639), .Y(n2406) );
  OAI21X1 U596 ( .A(n10758), .B(n10810), .C(n5757), .Y(n2407) );
  OAI21X1 U598 ( .A(n10758), .B(n10809), .C(n4958), .Y(n2408) );
  OAI21X1 U600 ( .A(n10758), .B(n10808), .C(n5067), .Y(n2409) );
  OAI21X1 U602 ( .A(n10757), .B(n10807), .C(n5176), .Y(n2410) );
  OAI21X1 U604 ( .A(n10757), .B(n10806), .C(n4535), .Y(n2411) );
  OAI21X1 U606 ( .A(n10757), .B(n10805), .C(n5756), .Y(n2412) );
  OAI21X1 U608 ( .A(n10757), .B(n10804), .C(n6022), .Y(n2413) );
  OAI21X1 U610 ( .A(n10757), .B(n10803), .C(n6154), .Y(n2414) );
  OAI21X1 U612 ( .A(n10758), .B(n10802), .C(n6286), .Y(n2415) );
  OAI21X1 U614 ( .A(n10757), .B(n10801), .C(n5402), .Y(n2416) );
  OAI21X1 U616 ( .A(n10758), .B(n10800), .C(n5520), .Y(n2417) );
  OAI21X1 U618 ( .A(n10757), .B(n10799), .C(n5638), .Y(n2418) );
  OAI21X1 U620 ( .A(n10757), .B(n10798), .C(n5890), .Y(n2419) );
  OAI21X1 U622 ( .A(n10757), .B(n10797), .C(n4957), .Y(n2420) );
  OAI21X1 U624 ( .A(n10758), .B(n10796), .C(n5066), .Y(n2421) );
  OAI21X1 U626 ( .A(n10757), .B(n10795), .C(n5175), .Y(n2422) );
  OAI21X1 U628 ( .A(n10757), .B(n10794), .C(n5285), .Y(n2423) );
  OAI21X1 U630 ( .A(n10758), .B(n10793), .C(n6021), .Y(n2424) );
  OAI21X1 U632 ( .A(n10757), .B(n10792), .C(n5519), .Y(n2425) );
  OAI21X1 U634 ( .A(n10757), .B(n10791), .C(n6153), .Y(n2426) );
  OAI21X1 U636 ( .A(n10757), .B(n10790), .C(n6285), .Y(n2427) );
  OAI21X1 U638 ( .A(n10758), .B(n10789), .C(n5401), .Y(n2428) );
  OAI21X1 U640 ( .A(n10758), .B(n10788), .C(n5284), .Y(n2429) );
  OAI21X1 U642 ( .A(n10757), .B(n10787), .C(n5637), .Y(n2430) );
  OAI21X1 U644 ( .A(n10758), .B(n10786), .C(n4956), .Y(n2431) );
  OAI21X1 U646 ( .A(n10758), .B(n10785), .C(n5889), .Y(n2432) );
  OAI21X1 U648 ( .A(n10757), .B(n10784), .C(n4534), .Y(n2433) );
  OAI21X1 U650 ( .A(n10757), .B(n10783), .C(n5755), .Y(n2434) );
  OAI21X1 U652 ( .A(n10757), .B(n10782), .C(n4641), .Y(n2435) );
  OAI21X1 U654 ( .A(n10758), .B(n10781), .C(n4749), .Y(n2436) );
  OAI21X1 U656 ( .A(n10758), .B(n10780), .C(n4854), .Y(n2437) );
  OAI21X1 U658 ( .A(n10757), .B(n10779), .C(n4416), .Y(n2438) );
  OAI21X1 U660 ( .A(n10758), .B(n10778), .C(n4415), .Y(n2439) );
  OAI21X1 U662 ( .A(n10758), .B(n10777), .C(n4748), .Y(n2440) );
  OAI21X1 U664 ( .A(n10757), .B(n10776), .C(n4414), .Y(n2441) );
  OAI21X1 U666 ( .A(n10758), .B(n10775), .C(n4413), .Y(n2442) );
  OAI21X1 U668 ( .A(n10758), .B(n10774), .C(n5174), .Y(n2443) );
  OAI21X1 U670 ( .A(n10757), .B(n10773), .C(n4533), .Y(n2444) );
  OAI21X1 U672 ( .A(n10758), .B(n10772), .C(n4640), .Y(n2445) );
  OAI21X1 U674 ( .A(n10757), .B(n10771), .C(n5283), .Y(n2446) );
  OAI21X1 U676 ( .A(n10757), .B(n10770), .C(n4412), .Y(n2447) );
  OAI21X1 U678 ( .A(n10757), .B(n10769), .C(n4747), .Y(n2448) );
  OAI21X1 U680 ( .A(n10758), .B(n10768), .C(n4411), .Y(n2449) );
  OAI21X1 U682 ( .A(n10758), .B(n10767), .C(n5065), .Y(n2450) );
  OAI21X1 U684 ( .A(n5906), .B(n5653), .C(reset_n), .Y(n365) );
  OAI21X1 U685 ( .A(n10755), .B(n10830), .C(n5754), .Y(n2451) );
  OAI21X1 U687 ( .A(n10755), .B(n10829), .C(n5753), .Y(n2452) );
  OAI21X1 U689 ( .A(n10755), .B(n10828), .C(n5636), .Y(n2453) );
  OAI21X1 U691 ( .A(n10755), .B(n10827), .C(n5518), .Y(n2454) );
  OAI21X1 U693 ( .A(n10755), .B(n10826), .C(n5400), .Y(n2455) );
  OAI21X1 U695 ( .A(n10755), .B(n10825), .C(n6284), .Y(n2456) );
  OAI21X1 U697 ( .A(n10755), .B(n10824), .C(n6152), .Y(n2457) );
  OAI21X1 U699 ( .A(n10755), .B(n10823), .C(n6020), .Y(n2458) );
  OAI21X1 U701 ( .A(n10755), .B(n10822), .C(n5888), .Y(n2459) );
  OAI21X1 U703 ( .A(n10755), .B(n10821), .C(n4853), .Y(n2460) );
  OAI21X1 U705 ( .A(n10755), .B(n10820), .C(n4746), .Y(n2461) );
  OAI21X1 U707 ( .A(n10755), .B(n10819), .C(n4639), .Y(n2462) );
  OAI21X1 U709 ( .A(n10755), .B(n10818), .C(n4532), .Y(n2463) );
  OAI21X1 U711 ( .A(n10755), .B(n10817), .C(n5752), .Y(n2464) );
  OAI21X1 U713 ( .A(n10755), .B(n10816), .C(n5635), .Y(n2465) );
  OAI21X1 U715 ( .A(n10755), .B(n10815), .C(n5517), .Y(n2466) );
  OAI21X1 U717 ( .A(n10756), .B(n10814), .C(n5399), .Y(n2467) );
  OAI21X1 U719 ( .A(n10756), .B(n10813), .C(n6283), .Y(n2468) );
  OAI21X1 U721 ( .A(n10755), .B(n10812), .C(n6151), .Y(n2469) );
  OAI21X1 U723 ( .A(n10756), .B(n10811), .C(n6019), .Y(n2470) );
  OAI21X1 U725 ( .A(n10756), .B(n10810), .C(n5887), .Y(n2471) );
  OAI21X1 U727 ( .A(n10756), .B(n10809), .C(n4852), .Y(n2472) );
  OAI21X1 U729 ( .A(n10756), .B(n10808), .C(n4745), .Y(n2473) );
  OAI21X1 U731 ( .A(n10755), .B(n10807), .C(n4638), .Y(n2474) );
  OAI21X1 U733 ( .A(n10755), .B(n10806), .C(n5282), .Y(n2475) );
  OAI21X1 U735 ( .A(n10755), .B(n10805), .C(n5886), .Y(n2476) );
  OAI21X1 U737 ( .A(n10755), .B(n10804), .C(n5634), .Y(n2477) );
  OAI21X1 U739 ( .A(n10755), .B(n10803), .C(n5516), .Y(n2478) );
  OAI21X1 U741 ( .A(n10756), .B(n10802), .C(n5398), .Y(n2479) );
  OAI21X1 U743 ( .A(n10755), .B(n10801), .C(n6282), .Y(n2480) );
  OAI21X1 U745 ( .A(n10756), .B(n10800), .C(n6150), .Y(n2481) );
  OAI21X1 U747 ( .A(n10755), .B(n10799), .C(n6018), .Y(n2482) );
  OAI21X1 U749 ( .A(n10755), .B(n10798), .C(n5751), .Y(n2483) );
  OAI21X1 U751 ( .A(n10755), .B(n10797), .C(n4851), .Y(n2484) );
  OAI21X1 U753 ( .A(n10756), .B(n10796), .C(n4744), .Y(n2485) );
  OAI21X1 U755 ( .A(n10755), .B(n10795), .C(n4637), .Y(n2486) );
  OAI21X1 U757 ( .A(n10755), .B(n10794), .C(n4531), .Y(n2487) );
  OAI21X1 U759 ( .A(n10756), .B(n10793), .C(n5633), .Y(n2488) );
  OAI21X1 U761 ( .A(n10755), .B(n10792), .C(n6149), .Y(n2489) );
  OAI21X1 U763 ( .A(n10755), .B(n10791), .C(n5515), .Y(n2490) );
  OAI21X1 U765 ( .A(n10755), .B(n10790), .C(n5397), .Y(n2491) );
  OAI21X1 U767 ( .A(n10756), .B(n10789), .C(n6281), .Y(n2492) );
  OAI21X1 U769 ( .A(n10756), .B(n10788), .C(n4530), .Y(n2493) );
  OAI21X1 U771 ( .A(n10755), .B(n10787), .C(n6017), .Y(n2494) );
  OAI21X1 U773 ( .A(n10756), .B(n10786), .C(n4850), .Y(n2495) );
  OAI21X1 U775 ( .A(n10756), .B(n10785), .C(n5750), .Y(n2496) );
  OAI21X1 U777 ( .A(n10755), .B(n10784), .C(n5281), .Y(n2497) );
  OAI21X1 U779 ( .A(n10755), .B(n10783), .C(n5885), .Y(n2498) );
  OAI21X1 U781 ( .A(n10755), .B(n10782), .C(n5173), .Y(n2499) );
  OAI21X1 U783 ( .A(n10756), .B(n10781), .C(n5064), .Y(n2500) );
  OAI21X1 U785 ( .A(n10756), .B(n10780), .C(n4955), .Y(n2501) );
  OAI21X1 U787 ( .A(n10755), .B(n10779), .C(n4410), .Y(n2502) );
  OAI21X1 U789 ( .A(n10756), .B(n10778), .C(n4409), .Y(n2503) );
  OAI21X1 U791 ( .A(n10756), .B(n10777), .C(n5063), .Y(n2504) );
  OAI21X1 U793 ( .A(n10755), .B(n10776), .C(n4408), .Y(n2505) );
  OAI21X1 U795 ( .A(n10756), .B(n10775), .C(n4407), .Y(n2506) );
  OAI21X1 U797 ( .A(n10756), .B(n10774), .C(n4636), .Y(n2507) );
  OAI21X1 U799 ( .A(n10755), .B(n10773), .C(n5280), .Y(n2508) );
  OAI21X1 U801 ( .A(n10756), .B(n10772), .C(n5172), .Y(n2509) );
  OAI21X1 U803 ( .A(n10755), .B(n10771), .C(n4529), .Y(n2510) );
  OAI21X1 U805 ( .A(n10755), .B(n10770), .C(n4406), .Y(n2511) );
  OAI21X1 U807 ( .A(n10755), .B(n10769), .C(n5062), .Y(n2512) );
  OAI21X1 U809 ( .A(n10756), .B(n10768), .C(n4405), .Y(n2513) );
  OAI21X1 U811 ( .A(n10756), .B(n10767), .C(n4743), .Y(n2514) );
  OAI21X1 U813 ( .A(n5906), .B(n5771), .C(reset_n), .Y(n431) );
  OAI21X1 U814 ( .A(n10753), .B(n10830), .C(n5632), .Y(n2515) );
  OAI21X1 U816 ( .A(n10753), .B(n10829), .C(n5631), .Y(n2516) );
  OAI21X1 U818 ( .A(n10753), .B(n10828), .C(n5749), .Y(n2517) );
  OAI21X1 U820 ( .A(n10753), .B(n10827), .C(n5396), .Y(n2518) );
  OAI21X1 U822 ( .A(n10753), .B(n10826), .C(n5514), .Y(n2519) );
  OAI21X1 U824 ( .A(n10753), .B(n10825), .C(n6148), .Y(n2520) );
  OAI21X1 U826 ( .A(n10753), .B(n10824), .C(n6280), .Y(n2521) );
  OAI21X1 U828 ( .A(n10753), .B(n10823), .C(n5884), .Y(n2522) );
  OAI21X1 U830 ( .A(n10753), .B(n10822), .C(n6016), .Y(n2523) );
  OAI21X1 U832 ( .A(n10753), .B(n10821), .C(n4742), .Y(n2524) );
  OAI21X1 U834 ( .A(n10753), .B(n10820), .C(n4849), .Y(n2525) );
  OAI21X1 U836 ( .A(n10753), .B(n10819), .C(n4528), .Y(n2526) );
  OAI21X1 U838 ( .A(n10753), .B(n10818), .C(n4635), .Y(n2527) );
  OAI21X1 U840 ( .A(n10753), .B(n10817), .C(n5630), .Y(n2528) );
  OAI21X1 U842 ( .A(n10753), .B(n10816), .C(n5748), .Y(n2529) );
  OAI21X1 U844 ( .A(n10753), .B(n10815), .C(n5395), .Y(n2530) );
  OAI21X1 U846 ( .A(n10754), .B(n10814), .C(n5513), .Y(n2531) );
  OAI21X1 U848 ( .A(n10754), .B(n10813), .C(n6147), .Y(n2532) );
  OAI21X1 U850 ( .A(n10753), .B(n10812), .C(n6279), .Y(n2533) );
  OAI21X1 U852 ( .A(n10754), .B(n10811), .C(n5883), .Y(n2534) );
  OAI21X1 U854 ( .A(n10754), .B(n10810), .C(n6015), .Y(n2535) );
  OAI21X1 U856 ( .A(n10754), .B(n10809), .C(n4741), .Y(n2536) );
  OAI21X1 U858 ( .A(n10754), .B(n10808), .C(n4848), .Y(n2537) );
  OAI21X1 U860 ( .A(n10753), .B(n10807), .C(n4527), .Y(n2538) );
  OAI21X1 U862 ( .A(n10753), .B(n10806), .C(n5171), .Y(n2539) );
  OAI21X1 U864 ( .A(n10753), .B(n10805), .C(n6014), .Y(n2540) );
  OAI21X1 U866 ( .A(n10753), .B(n10804), .C(n5747), .Y(n2541) );
  OAI21X1 U868 ( .A(n10753), .B(n10803), .C(n5394), .Y(n2542) );
  OAI21X1 U870 ( .A(n10754), .B(n10802), .C(n5512), .Y(n2543) );
  OAI21X1 U872 ( .A(n10753), .B(n10801), .C(n6146), .Y(n2544) );
  OAI21X1 U874 ( .A(n10754), .B(n10800), .C(n6278), .Y(n2545) );
  OAI21X1 U876 ( .A(n10753), .B(n10799), .C(n5882), .Y(n2546) );
  OAI21X1 U878 ( .A(n10753), .B(n10798), .C(n5629), .Y(n2547) );
  OAI21X1 U880 ( .A(n10753), .B(n10797), .C(n4740), .Y(n2548) );
  OAI21X1 U882 ( .A(n10754), .B(n10796), .C(n4847), .Y(n2549) );
  OAI21X1 U884 ( .A(n10753), .B(n10795), .C(n4526), .Y(n2550) );
  OAI21X1 U886 ( .A(n10753), .B(n10794), .C(n4634), .Y(n2551) );
  OAI21X1 U888 ( .A(n10754), .B(n10793), .C(n5746), .Y(n2552) );
  OAI21X1 U890 ( .A(n10753), .B(n10792), .C(n6277), .Y(n2553) );
  OAI21X1 U892 ( .A(n10753), .B(n10791), .C(n5393), .Y(n2554) );
  OAI21X1 U894 ( .A(n10753), .B(n10790), .C(n5511), .Y(n2555) );
  OAI21X1 U896 ( .A(n10754), .B(n10789), .C(n6145), .Y(n2556) );
  OAI21X1 U898 ( .A(n10754), .B(n10788), .C(n4633), .Y(n2557) );
  OAI21X1 U900 ( .A(n10753), .B(n10787), .C(n5881), .Y(n2558) );
  OAI21X1 U902 ( .A(n10754), .B(n10786), .C(n4739), .Y(n2559) );
  OAI21X1 U904 ( .A(n10754), .B(n10785), .C(n5628), .Y(n2560) );
  OAI21X1 U906 ( .A(n10753), .B(n10784), .C(n5170), .Y(n2561) );
  OAI21X1 U908 ( .A(n10753), .B(n10783), .C(n6013), .Y(n2562) );
  OAI21X1 U910 ( .A(n10753), .B(n10782), .C(n5279), .Y(n2563) );
  OAI21X1 U912 ( .A(n10754), .B(n10781), .C(n4954), .Y(n2564) );
  OAI21X1 U914 ( .A(n10754), .B(n10780), .C(n5061), .Y(n2565) );
  OAI21X1 U916 ( .A(n10753), .B(n10779), .C(n4404), .Y(n2566) );
  OAI21X1 U918 ( .A(n10754), .B(n10778), .C(n4403), .Y(n2567) );
  OAI21X1 U920 ( .A(n10754), .B(n10777), .C(n4953), .Y(n2568) );
  OAI21X1 U922 ( .A(n10753), .B(n10776), .C(n4402), .Y(n2569) );
  OAI21X1 U924 ( .A(n10754), .B(n10775), .C(n4401), .Y(n2570) );
  OAI21X1 U926 ( .A(n10754), .B(n10774), .C(n4525), .Y(n2571) );
  OAI21X1 U928 ( .A(n10753), .B(n10773), .C(n5169), .Y(n2572) );
  OAI21X1 U930 ( .A(n10754), .B(n10772), .C(n5278), .Y(n2573) );
  OAI21X1 U932 ( .A(n10753), .B(n10771), .C(n4632), .Y(n2574) );
  OAI21X1 U934 ( .A(n10753), .B(n10770), .C(n4400), .Y(n2575) );
  OAI21X1 U936 ( .A(n10753), .B(n10769), .C(n4952), .Y(n2576) );
  OAI21X1 U938 ( .A(n10754), .B(n10768), .C(n4399), .Y(n2577) );
  OAI21X1 U940 ( .A(n10754), .B(n10767), .C(n4846), .Y(n2578) );
  OAI21X1 U942 ( .A(n5906), .B(n5535), .C(reset_n), .Y(n497) );
  OAI21X1 U943 ( .A(n10751), .B(n10830), .C(n5510), .Y(n2579) );
  OAI21X1 U945 ( .A(n10751), .B(n10829), .C(n5509), .Y(n2580) );
  OAI21X1 U947 ( .A(n10751), .B(n10828), .C(n5392), .Y(n2581) );
  OAI21X1 U949 ( .A(n10751), .B(n10827), .C(n5745), .Y(n2582) );
  OAI21X1 U951 ( .A(n10751), .B(n10826), .C(n5627), .Y(n2583) );
  OAI21X1 U953 ( .A(n10751), .B(n10825), .C(n6012), .Y(n2584) );
  OAI21X1 U955 ( .A(n10751), .B(n10824), .C(n5880), .Y(n2585) );
  OAI21X1 U957 ( .A(n10751), .B(n10823), .C(n6276), .Y(n2586) );
  OAI21X1 U959 ( .A(n10751), .B(n10822), .C(n6144), .Y(n2587) );
  OAI21X1 U961 ( .A(n10751), .B(n10821), .C(n4631), .Y(n2588) );
  OAI21X1 U963 ( .A(n10751), .B(n10820), .C(n4524), .Y(n2589) );
  OAI21X1 U965 ( .A(n10751), .B(n10819), .C(n4845), .Y(n2590) );
  OAI21X1 U967 ( .A(n10751), .B(n10818), .C(n4738), .Y(n2591) );
  OAI21X1 U969 ( .A(n10751), .B(n10817), .C(n5508), .Y(n2592) );
  OAI21X1 U971 ( .A(n10751), .B(n10816), .C(n5391), .Y(n2593) );
  OAI21X1 U973 ( .A(n10751), .B(n10815), .C(n5744), .Y(n2594) );
  OAI21X1 U975 ( .A(n10752), .B(n10814), .C(n5626), .Y(n2595) );
  OAI21X1 U977 ( .A(n10752), .B(n10813), .C(n6011), .Y(n2596) );
  OAI21X1 U979 ( .A(n10751), .B(n10812), .C(n5879), .Y(n2597) );
  OAI21X1 U981 ( .A(n10752), .B(n10811), .C(n6275), .Y(n2598) );
  OAI21X1 U983 ( .A(n10752), .B(n10810), .C(n6143), .Y(n2599) );
  OAI21X1 U985 ( .A(n10752), .B(n10809), .C(n4630), .Y(n2600) );
  OAI21X1 U987 ( .A(n10752), .B(n10808), .C(n4523), .Y(n2601) );
  OAI21X1 U989 ( .A(n10751), .B(n10807), .C(n4844), .Y(n2602) );
  OAI21X1 U991 ( .A(n10751), .B(n10806), .C(n5060), .Y(n2603) );
  OAI21X1 U993 ( .A(n10751), .B(n10805), .C(n6142), .Y(n2604) );
  OAI21X1 U995 ( .A(n10751), .B(n10804), .C(n5390), .Y(n2605) );
  OAI21X1 U997 ( .A(n10751), .B(n10803), .C(n5743), .Y(n2606) );
  OAI21X1 U999 ( .A(n10752), .B(n10802), .C(n5625), .Y(n2607) );
  OAI21X1 U1001 ( .A(n10751), .B(n10801), .C(n6010), .Y(n2608) );
  OAI21X1 U1003 ( .A(n10752), .B(n10800), .C(n5878), .Y(n2609) );
  OAI21X1 U1005 ( .A(n10751), .B(n10799), .C(n6274), .Y(n2610) );
  OAI21X1 U1007 ( .A(n10751), .B(n10798), .C(n5507), .Y(n2611) );
  OAI21X1 U1009 ( .A(n10751), .B(n10797), .C(n4629), .Y(n2612) );
  OAI21X1 U1011 ( .A(n10752), .B(n10796), .C(n4522), .Y(n2613) );
  OAI21X1 U1013 ( .A(n10751), .B(n10795), .C(n4843), .Y(n2614) );
  OAI21X1 U1015 ( .A(n10751), .B(n10794), .C(n4737), .Y(n2615) );
  OAI21X1 U1017 ( .A(n10752), .B(n10793), .C(n5389), .Y(n2616) );
  OAI21X1 U1019 ( .A(n10751), .B(n10792), .C(n5877), .Y(n2617) );
  OAI21X1 U1021 ( .A(n10751), .B(n10791), .C(n5742), .Y(n2618) );
  OAI21X1 U1023 ( .A(n10751), .B(n10790), .C(n5624), .Y(n2619) );
  OAI21X1 U1025 ( .A(n10752), .B(n10789), .C(n6009), .Y(n2620) );
  OAI21X1 U1027 ( .A(n10752), .B(n10788), .C(n4736), .Y(n2621) );
  OAI21X1 U1029 ( .A(n10751), .B(n10787), .C(n6273), .Y(n2622) );
  OAI21X1 U1031 ( .A(n10752), .B(n10786), .C(n4628), .Y(n2623) );
  OAI21X1 U1033 ( .A(n10752), .B(n10785), .C(n5506), .Y(n2624) );
  OAI21X1 U1035 ( .A(n10751), .B(n10784), .C(n5059), .Y(n2625) );
  OAI21X1 U1037 ( .A(n10751), .B(n10783), .C(n6141), .Y(n2626) );
  OAI21X1 U1039 ( .A(n10751), .B(n10782), .C(n4951), .Y(n2627) );
  OAI21X1 U1041 ( .A(n10752), .B(n10781), .C(n5277), .Y(n2628) );
  OAI21X1 U1043 ( .A(n10752), .B(n10780), .C(n5168), .Y(n2629) );
  OAI21X1 U1045 ( .A(n10751), .B(n10779), .C(n4398), .Y(n2630) );
  OAI21X1 U1047 ( .A(n10752), .B(n10778), .C(n4397), .Y(n2631) );
  OAI21X1 U1049 ( .A(n10752), .B(n10777), .C(n5276), .Y(n2632) );
  OAI21X1 U1051 ( .A(n10751), .B(n10776), .C(n4396), .Y(n2633) );
  OAI21X1 U1053 ( .A(n10752), .B(n10775), .C(n4395), .Y(n2634) );
  OAI21X1 U1055 ( .A(n10752), .B(n10774), .C(n4842), .Y(n2635) );
  OAI21X1 U1057 ( .A(n10751), .B(n10773), .C(n5058), .Y(n2636) );
  OAI21X1 U1059 ( .A(n10752), .B(n10772), .C(n4950), .Y(n2637) );
  OAI21X1 U1061 ( .A(n10751), .B(n10771), .C(n4735), .Y(n2638) );
  OAI21X1 U1063 ( .A(n10751), .B(n10770), .C(n4394), .Y(n2639) );
  OAI21X1 U1065 ( .A(n10751), .B(n10769), .C(n5275), .Y(n2640) );
  OAI21X1 U1067 ( .A(n10752), .B(n10768), .C(n4393), .Y(n2641) );
  OAI21X1 U1069 ( .A(n10752), .B(n10767), .C(n4521), .Y(n2642) );
  OAI21X1 U1071 ( .A(n5906), .B(n5417), .C(reset_n), .Y(n563) );
  OAI21X1 U1072 ( .A(n10749), .B(n10830), .C(n5388), .Y(n2643) );
  OAI21X1 U1074 ( .A(n10749), .B(n10829), .C(n5387), .Y(n2644) );
  OAI21X1 U1076 ( .A(n10749), .B(n10828), .C(n5505), .Y(n2645) );
  OAI21X1 U1078 ( .A(n10749), .B(n10827), .C(n5623), .Y(n2646) );
  OAI21X1 U1080 ( .A(n10749), .B(n10826), .C(n5741), .Y(n2647) );
  OAI21X1 U1082 ( .A(n10749), .B(n10825), .C(n5876), .Y(n2648) );
  OAI21X1 U1084 ( .A(n10749), .B(n10824), .C(n6008), .Y(n2649) );
  OAI21X1 U1086 ( .A(n10749), .B(n10823), .C(n6140), .Y(n2650) );
  OAI21X1 U1088 ( .A(n10749), .B(n10822), .C(n6272), .Y(n2651) );
  OAI21X1 U1090 ( .A(n10749), .B(n10821), .C(n4520), .Y(n2652) );
  OAI21X1 U1092 ( .A(n10749), .B(n10820), .C(n4627), .Y(n2653) );
  OAI21X1 U1094 ( .A(n10749), .B(n10819), .C(n4734), .Y(n2654) );
  OAI21X1 U1096 ( .A(n10749), .B(n10818), .C(n4841), .Y(n2655) );
  OAI21X1 U1098 ( .A(n10749), .B(n10817), .C(n5386), .Y(n2656) );
  OAI21X1 U1100 ( .A(n10749), .B(n10816), .C(n5504), .Y(n2657) );
  OAI21X1 U1102 ( .A(n10750), .B(n10815), .C(n5622), .Y(n2658) );
  OAI21X1 U1104 ( .A(n10749), .B(n10814), .C(n5740), .Y(n2659) );
  OAI21X1 U1106 ( .A(n10750), .B(n10813), .C(n5875), .Y(n2660) );
  OAI21X1 U1108 ( .A(n10749), .B(n10812), .C(n6007), .Y(n2661) );
  OAI21X1 U1110 ( .A(n10750), .B(n10811), .C(n6139), .Y(n2662) );
  OAI21X1 U1112 ( .A(n10750), .B(n10810), .C(n6271), .Y(n2663) );
  OAI21X1 U1114 ( .A(n10750), .B(n10809), .C(n4519), .Y(n2664) );
  OAI21X1 U1116 ( .A(n10750), .B(n10808), .C(n4626), .Y(n2665) );
  OAI21X1 U1118 ( .A(n10749), .B(n10807), .C(n4733), .Y(n2666) );
  OAI21X1 U1120 ( .A(n10749), .B(n10806), .C(n4949), .Y(n2667) );
  OAI21X1 U1122 ( .A(n10749), .B(n10805), .C(n6270), .Y(n2668) );
  OAI21X1 U1124 ( .A(n10749), .B(n10804), .C(n5503), .Y(n2669) );
  OAI21X1 U1126 ( .A(n10749), .B(n10803), .C(n5621), .Y(n2670) );
  OAI21X1 U1128 ( .A(n10750), .B(n10802), .C(n5739), .Y(n2671) );
  OAI21X1 U1130 ( .A(n10750), .B(n10801), .C(n5874), .Y(n2672) );
  OAI21X1 U1132 ( .A(n10750), .B(n10800), .C(n6006), .Y(n2673) );
  OAI21X1 U1134 ( .A(n10749), .B(n10799), .C(n6138), .Y(n2674) );
  OAI21X1 U1136 ( .A(n10749), .B(n10798), .C(n5385), .Y(n2675) );
  OAI21X1 U1138 ( .A(n10749), .B(n10797), .C(n4518), .Y(n2676) );
  OAI21X1 U1140 ( .A(n10749), .B(n10796), .C(n4625), .Y(n2677) );
  OAI21X1 U1142 ( .A(n10750), .B(n10795), .C(n4732), .Y(n2678) );
  OAI21X1 U1144 ( .A(n10749), .B(n10794), .C(n4840), .Y(n2679) );
  OAI21X1 U1146 ( .A(n10749), .B(n10793), .C(n5502), .Y(n2680) );
  OAI21X1 U1148 ( .A(n10749), .B(n10792), .C(n6005), .Y(n2681) );
  OAI21X1 U1150 ( .A(n10749), .B(n10791), .C(n5620), .Y(n2682) );
  OAI21X1 U1152 ( .A(n10749), .B(n10790), .C(n5738), .Y(n2683) );
  OAI21X1 U1154 ( .A(n10750), .B(n10789), .C(n5873), .Y(n2684) );
  OAI21X1 U1156 ( .A(n10750), .B(n10788), .C(n4839), .Y(n2685) );
  OAI21X1 U1158 ( .A(n10749), .B(n10787), .C(n6137), .Y(n2686) );
  OAI21X1 U1160 ( .A(n10750), .B(n10786), .C(n4517), .Y(n2687) );
  OAI21X1 U1162 ( .A(n10750), .B(n10785), .C(n5384), .Y(n2688) );
  OAI21X1 U1164 ( .A(n10749), .B(n10784), .C(n4948), .Y(n2689) );
  OAI21X1 U1166 ( .A(n10750), .B(n10783), .C(n6269), .Y(n2690) );
  OAI21X1 U1168 ( .A(n10749), .B(n10782), .C(n5057), .Y(n2691) );
  OAI21X1 U1170 ( .A(n10750), .B(n10781), .C(n5167), .Y(n2692) );
  OAI21X1 U1172 ( .A(n10750), .B(n10780), .C(n5274), .Y(n2693) );
  OAI21X1 U1174 ( .A(n10750), .B(n10779), .C(n4392), .Y(n2694) );
  OAI21X1 U1176 ( .A(n10749), .B(n10778), .C(n4391), .Y(n2695) );
  OAI21X1 U1178 ( .A(n10749), .B(n10777), .C(n5166), .Y(n2696) );
  OAI21X1 U1180 ( .A(n10749), .B(n10776), .C(n4390), .Y(n2697) );
  OAI21X1 U1182 ( .A(n10750), .B(n10775), .C(n4389), .Y(n2698) );
  OAI21X1 U1184 ( .A(n10750), .B(n10774), .C(n4731), .Y(n2699) );
  OAI21X1 U1186 ( .A(n10749), .B(n10773), .C(n4947), .Y(n2700) );
  OAI21X1 U1188 ( .A(n10750), .B(n10772), .C(n5056), .Y(n2701) );
  OAI21X1 U1190 ( .A(n10749), .B(n10771), .C(n4838), .Y(n2702) );
  OAI21X1 U1192 ( .A(n10749), .B(n10770), .C(n4388), .Y(n2703) );
  OAI21X1 U1194 ( .A(n10749), .B(n10769), .C(n5165), .Y(n2704) );
  OAI21X1 U1196 ( .A(n10750), .B(n10768), .C(n4387), .Y(n2705) );
  OAI21X1 U1198 ( .A(n10750), .B(n10767), .C(n4624), .Y(n2706) );
  OAI21X1 U1200 ( .A(n5906), .B(n5299), .C(reset_n), .Y(n629) );
  NAND3X1 U1201 ( .A(waddr[3]), .B(n631), .C(waddr[4]), .Y(n167) );
  OAI21X1 U1202 ( .A(n10747), .B(n10830), .C(n6268), .Y(n2707) );
  OAI21X1 U1204 ( .A(n10747), .B(n10829), .C(n6267), .Y(n2708) );
  OAI21X1 U1206 ( .A(n10747), .B(n10828), .C(n6136), .Y(n2709) );
  OAI21X1 U1208 ( .A(n10747), .B(n10827), .C(n6004), .Y(n2710) );
  OAI21X1 U1210 ( .A(n10747), .B(n10826), .C(n5872), .Y(n2711) );
  OAI21X1 U1212 ( .A(n10747), .B(n10825), .C(n5737), .Y(n2712) );
  OAI21X1 U1214 ( .A(n10747), .B(n10824), .C(n5619), .Y(n2713) );
  OAI21X1 U1216 ( .A(n10747), .B(n10823), .C(n5501), .Y(n2714) );
  OAI21X1 U1218 ( .A(n10747), .B(n10822), .C(n5383), .Y(n2715) );
  OAI21X1 U1220 ( .A(n10747), .B(n10821), .C(n5273), .Y(n2716) );
  OAI21X1 U1222 ( .A(n10747), .B(n10820), .C(n5164), .Y(n2717) );
  OAI21X1 U1224 ( .A(n10747), .B(n10819), .C(n5055), .Y(n2718) );
  OAI21X1 U1226 ( .A(n10747), .B(n10818), .C(n4946), .Y(n2719) );
  OAI21X1 U1228 ( .A(n10747), .B(n10817), .C(n6266), .Y(n2720) );
  OAI21X1 U1230 ( .A(n10747), .B(n10816), .C(n6135), .Y(n2721) );
  OAI21X1 U1232 ( .A(n10747), .B(n10815), .C(n6003), .Y(n2722) );
  OAI21X1 U1234 ( .A(n10748), .B(n10814), .C(n5871), .Y(n2723) );
  OAI21X1 U1236 ( .A(n10748), .B(n10813), .C(n5736), .Y(n2724) );
  OAI21X1 U1238 ( .A(n10747), .B(n10812), .C(n5618), .Y(n2725) );
  OAI21X1 U1240 ( .A(n10748), .B(n10811), .C(n5500), .Y(n2726) );
  OAI21X1 U1242 ( .A(n10748), .B(n10810), .C(n5382), .Y(n2727) );
  OAI21X1 U1244 ( .A(n10748), .B(n10809), .C(n5272), .Y(n2728) );
  OAI21X1 U1246 ( .A(n10748), .B(n10808), .C(n5163), .Y(n2729) );
  OAI21X1 U1248 ( .A(n10747), .B(n10807), .C(n5054), .Y(n2730) );
  OAI21X1 U1250 ( .A(n10747), .B(n10806), .C(n4837), .Y(n2731) );
  OAI21X1 U1252 ( .A(n10747), .B(n10805), .C(n5381), .Y(n2732) );
  OAI21X1 U1254 ( .A(n10747), .B(n10804), .C(n6134), .Y(n2733) );
  OAI21X1 U1256 ( .A(n10747), .B(n10803), .C(n6002), .Y(n2734) );
  OAI21X1 U1258 ( .A(n10748), .B(n10802), .C(n5870), .Y(n2735) );
  OAI21X1 U1260 ( .A(n10747), .B(n10801), .C(n5735), .Y(n2736) );
  OAI21X1 U1262 ( .A(n10748), .B(n10800), .C(n5617), .Y(n2737) );
  OAI21X1 U1264 ( .A(n10747), .B(n10799), .C(n5499), .Y(n2738) );
  OAI21X1 U1266 ( .A(n10747), .B(n10798), .C(n6265), .Y(n2739) );
  OAI21X1 U1268 ( .A(n10747), .B(n10797), .C(n5271), .Y(n2740) );
  OAI21X1 U1270 ( .A(n10748), .B(n10796), .C(n5162), .Y(n2741) );
  OAI21X1 U1272 ( .A(n10747), .B(n10795), .C(n5053), .Y(n2742) );
  OAI21X1 U1274 ( .A(n10747), .B(n10794), .C(n4945), .Y(n2743) );
  OAI21X1 U1276 ( .A(n10748), .B(n10793), .C(n6133), .Y(n2744) );
  OAI21X1 U1278 ( .A(n10747), .B(n10792), .C(n5616), .Y(n2745) );
  OAI21X1 U1280 ( .A(n10747), .B(n10791), .C(n6001), .Y(n2746) );
  OAI21X1 U1282 ( .A(n10747), .B(n10790), .C(n5869), .Y(n2747) );
  OAI21X1 U1284 ( .A(n10748), .B(n10789), .C(n5734), .Y(n2748) );
  OAI21X1 U1286 ( .A(n10748), .B(n10788), .C(n4944), .Y(n2749) );
  OAI21X1 U1288 ( .A(n10747), .B(n10787), .C(n5498), .Y(n2750) );
  OAI21X1 U1290 ( .A(n10748), .B(n10786), .C(n5270), .Y(n2751) );
  OAI21X1 U1292 ( .A(n10748), .B(n10785), .C(n6264), .Y(n2752) );
  OAI21X1 U1294 ( .A(n10747), .B(n10784), .C(n4836), .Y(n2753) );
  OAI21X1 U1296 ( .A(n10747), .B(n10783), .C(n5380), .Y(n2754) );
  OAI21X1 U1298 ( .A(n10747), .B(n10782), .C(n4730), .Y(n2755) );
  OAI21X1 U1300 ( .A(n10748), .B(n10781), .C(n4623), .Y(n2756) );
  OAI21X1 U1302 ( .A(n10748), .B(n10780), .C(n4516), .Y(n2757) );
  OAI21X1 U1304 ( .A(n10747), .B(n10779), .C(n4386), .Y(n2758) );
  OAI21X1 U1306 ( .A(n10748), .B(n10778), .C(n4385), .Y(n2759) );
  OAI21X1 U1308 ( .A(n10748), .B(n10777), .C(n4622), .Y(n2760) );
  OAI21X1 U1310 ( .A(n10747), .B(n10776), .C(n4384), .Y(n2761) );
  OAI21X1 U1312 ( .A(n10748), .B(n10775), .C(n4383), .Y(n2762) );
  OAI21X1 U1314 ( .A(n10748), .B(n10774), .C(n5052), .Y(n2763) );
  OAI21X1 U1316 ( .A(n10747), .B(n10773), .C(n4835), .Y(n2764) );
  OAI21X1 U1318 ( .A(n10748), .B(n10772), .C(n4729), .Y(n2765) );
  OAI21X1 U1320 ( .A(n10747), .B(n10771), .C(n4943), .Y(n2766) );
  OAI21X1 U1322 ( .A(n10747), .B(n10770), .C(n4382), .Y(n2767) );
  OAI21X1 U1324 ( .A(n10747), .B(n10769), .C(n4621), .Y(n2768) );
  OAI21X1 U1326 ( .A(n10748), .B(n10768), .C(n4381), .Y(n2769) );
  OAI21X1 U1328 ( .A(n10748), .B(n10767), .C(n5161), .Y(n2770) );
  OAI21X1 U1330 ( .A(n5774), .B(n6302), .C(reset_n), .Y(n696) );
  OAI21X1 U1331 ( .A(n10745), .B(n10830), .C(n6132), .Y(n2771) );
  OAI21X1 U1333 ( .A(n10745), .B(n10829), .C(n6131), .Y(n2772) );
  OAI21X1 U1335 ( .A(n10745), .B(n10828), .C(n6263), .Y(n2773) );
  OAI21X1 U1337 ( .A(n10745), .B(n10827), .C(n5868), .Y(n2774) );
  OAI21X1 U1339 ( .A(n10745), .B(n10826), .C(n6000), .Y(n2775) );
  OAI21X1 U1341 ( .A(n10745), .B(n10825), .C(n5615), .Y(n2776) );
  OAI21X1 U1343 ( .A(n10745), .B(n10824), .C(n5733), .Y(n2777) );
  OAI21X1 U1345 ( .A(n10745), .B(n10823), .C(n5379), .Y(n2778) );
  OAI21X1 U1347 ( .A(n10745), .B(n10822), .C(n5497), .Y(n2779) );
  OAI21X1 U1349 ( .A(n10745), .B(n10821), .C(n5160), .Y(n2780) );
  OAI21X1 U1351 ( .A(n10745), .B(n10820), .C(n5269), .Y(n2781) );
  OAI21X1 U1353 ( .A(n10745), .B(n10819), .C(n4942), .Y(n2782) );
  OAI21X1 U1355 ( .A(n10745), .B(n10818), .C(n5051), .Y(n2783) );
  OAI21X1 U1357 ( .A(n10745), .B(n10817), .C(n6130), .Y(n2784) );
  OAI21X1 U1359 ( .A(n10745), .B(n10816), .C(n6262), .Y(n2785) );
  OAI21X1 U1361 ( .A(n10745), .B(n10815), .C(n5867), .Y(n2786) );
  OAI21X1 U1363 ( .A(n10746), .B(n10814), .C(n5999), .Y(n2787) );
  OAI21X1 U1365 ( .A(n10746), .B(n10813), .C(n5614), .Y(n2788) );
  OAI21X1 U1367 ( .A(n10745), .B(n10812), .C(n5732), .Y(n2789) );
  OAI21X1 U1369 ( .A(n10746), .B(n10811), .C(n5378), .Y(n2790) );
  OAI21X1 U1371 ( .A(n10746), .B(n10810), .C(n5496), .Y(n2791) );
  OAI21X1 U1373 ( .A(n10746), .B(n10809), .C(n5159), .Y(n2792) );
  OAI21X1 U1375 ( .A(n10746), .B(n10808), .C(n5268), .Y(n2793) );
  OAI21X1 U1377 ( .A(n10745), .B(n10807), .C(n4941), .Y(n2794) );
  OAI21X1 U1379 ( .A(n10745), .B(n10806), .C(n4728), .Y(n2795) );
  OAI21X1 U1381 ( .A(n10745), .B(n10805), .C(n5495), .Y(n2796) );
  OAI21X1 U1383 ( .A(n10745), .B(n10804), .C(n6261), .Y(n2797) );
  OAI21X1 U1385 ( .A(n10745), .B(n10803), .C(n5866), .Y(n2798) );
  OAI21X1 U1387 ( .A(n10746), .B(n10802), .C(n5998), .Y(n2799) );
  OAI21X1 U1389 ( .A(n10745), .B(n10801), .C(n5613), .Y(n2800) );
  OAI21X1 U1391 ( .A(n10746), .B(n10800), .C(n5731), .Y(n2801) );
  OAI21X1 U1393 ( .A(n10745), .B(n10799), .C(n5377), .Y(n2802) );
  OAI21X1 U1395 ( .A(n10745), .B(n10798), .C(n6129), .Y(n2803) );
  OAI21X1 U1397 ( .A(n10745), .B(n10797), .C(n5158), .Y(n2804) );
  OAI21X1 U1399 ( .A(n10746), .B(n10796), .C(n5267), .Y(n2805) );
  OAI21X1 U1401 ( .A(n10745), .B(n10795), .C(n4940), .Y(n2806) );
  OAI21X1 U1403 ( .A(n10745), .B(n10794), .C(n5050), .Y(n2807) );
  OAI21X1 U1405 ( .A(n10746), .B(n10793), .C(n6260), .Y(n2808) );
  OAI21X1 U1407 ( .A(n10745), .B(n10792), .C(n5730), .Y(n2809) );
  OAI21X1 U1409 ( .A(n10745), .B(n10791), .C(n5865), .Y(n2810) );
  OAI21X1 U1411 ( .A(n10745), .B(n10790), .C(n5997), .Y(n2811) );
  OAI21X1 U1413 ( .A(n10746), .B(n10789), .C(n5612), .Y(n2812) );
  OAI21X1 U1415 ( .A(n10746), .B(n10788), .C(n5049), .Y(n2813) );
  OAI21X1 U1417 ( .A(n10745), .B(n10787), .C(n5376), .Y(n2814) );
  OAI21X1 U1419 ( .A(n10746), .B(n10786), .C(n5157), .Y(n2815) );
  OAI21X1 U1421 ( .A(n10746), .B(n10785), .C(n6128), .Y(n2816) );
  OAI21X1 U1423 ( .A(n10745), .B(n10784), .C(n4727), .Y(n2817) );
  OAI21X1 U1425 ( .A(n10745), .B(n10783), .C(n5494), .Y(n2818) );
  OAI21X1 U1427 ( .A(n10745), .B(n10782), .C(n4834), .Y(n2819) );
  OAI21X1 U1429 ( .A(n10746), .B(n10781), .C(n4515), .Y(n2820) );
  OAI21X1 U1431 ( .A(n10746), .B(n10780), .C(n4620), .Y(n2821) );
  OAI21X1 U1433 ( .A(n10745), .B(n10779), .C(n4380), .Y(n2822) );
  OAI21X1 U1435 ( .A(n10746), .B(n10778), .C(n4379), .Y(n2823) );
  OAI21X1 U1437 ( .A(n10746), .B(n10777), .C(n4514), .Y(n2824) );
  OAI21X1 U1439 ( .A(n10745), .B(n10776), .C(n4378), .Y(n2825) );
  OAI21X1 U1441 ( .A(n10746), .B(n10775), .C(n4377), .Y(n2826) );
  OAI21X1 U1443 ( .A(n10746), .B(n10774), .C(n4939), .Y(n2827) );
  OAI21X1 U1445 ( .A(n10745), .B(n10773), .C(n4726), .Y(n2828) );
  OAI21X1 U1447 ( .A(n10746), .B(n10772), .C(n4833), .Y(n2829) );
  OAI21X1 U1449 ( .A(n10745), .B(n10771), .C(n5048), .Y(n2830) );
  OAI21X1 U1451 ( .A(n10745), .B(n10770), .C(n4376), .Y(n2831) );
  OAI21X1 U1453 ( .A(n10745), .B(n10769), .C(n4513), .Y(n2832) );
  OAI21X1 U1455 ( .A(n10746), .B(n10768), .C(n4375), .Y(n2833) );
  OAI21X1 U1457 ( .A(n10746), .B(n10767), .C(n5266), .Y(n2834) );
  OAI21X1 U1459 ( .A(n5773), .B(n6302), .C(reset_n), .Y(n762) );
  OAI21X1 U1460 ( .A(n10743), .B(n10830), .C(n5996), .Y(n2835) );
  OAI21X1 U1462 ( .A(n10743), .B(n10829), .C(n5995), .Y(n2836) );
  OAI21X1 U1464 ( .A(n10743), .B(n10828), .C(n5864), .Y(n2837) );
  OAI21X1 U1466 ( .A(n10743), .B(n10827), .C(n6259), .Y(n2838) );
  OAI21X1 U1468 ( .A(n10743), .B(n10826), .C(n6127), .Y(n2839) );
  OAI21X1 U1470 ( .A(n10743), .B(n10825), .C(n5493), .Y(n2840) );
  OAI21X1 U1472 ( .A(n10743), .B(n10824), .C(n5375), .Y(n2841) );
  OAI21X1 U1474 ( .A(n10743), .B(n10823), .C(n5729), .Y(n2842) );
  OAI21X1 U1476 ( .A(n10743), .B(n10822), .C(n5611), .Y(n2843) );
  OAI21X1 U1478 ( .A(n10743), .B(n10821), .C(n5047), .Y(n2844) );
  OAI21X1 U1480 ( .A(n10743), .B(n10820), .C(n4938), .Y(n2845) );
  OAI21X1 U1482 ( .A(n10743), .B(n10819), .C(n5265), .Y(n2846) );
  OAI21X1 U1484 ( .A(n10743), .B(n10818), .C(n5156), .Y(n2847) );
  OAI21X1 U1486 ( .A(n10743), .B(n10817), .C(n5994), .Y(n2848) );
  OAI21X1 U1488 ( .A(n10743), .B(n10816), .C(n5863), .Y(n2849) );
  OAI21X1 U1490 ( .A(n10743), .B(n10815), .C(n6258), .Y(n2850) );
  OAI21X1 U1492 ( .A(n10744), .B(n10814), .C(n6126), .Y(n2851) );
  OAI21X1 U1494 ( .A(n10744), .B(n10813), .C(n5492), .Y(n2852) );
  OAI21X1 U1496 ( .A(n10743), .B(n10812), .C(n5374), .Y(n2853) );
  OAI21X1 U1498 ( .A(n10744), .B(n10811), .C(n5728), .Y(n2854) );
  OAI21X1 U1500 ( .A(n10744), .B(n10810), .C(n5610), .Y(n2855) );
  OAI21X1 U1502 ( .A(n10744), .B(n10809), .C(n5046), .Y(n2856) );
  OAI21X1 U1504 ( .A(n10744), .B(n10808), .C(n4937), .Y(n2857) );
  OAI21X1 U1506 ( .A(n10743), .B(n10807), .C(n5264), .Y(n2858) );
  OAI21X1 U1508 ( .A(n10743), .B(n10806), .C(n4619), .Y(n2859) );
  OAI21X1 U1510 ( .A(n10743), .B(n10805), .C(n5609), .Y(n2860) );
  OAI21X1 U1512 ( .A(n10743), .B(n10804), .C(n5862), .Y(n2861) );
  OAI21X1 U1514 ( .A(n10743), .B(n10803), .C(n6257), .Y(n2862) );
  OAI21X1 U1516 ( .A(n10744), .B(n10802), .C(n6125), .Y(n2863) );
  OAI21X1 U1518 ( .A(n10743), .B(n10801), .C(n5491), .Y(n2864) );
  OAI21X1 U1520 ( .A(n10744), .B(n10800), .C(n5373), .Y(n2865) );
  OAI21X1 U1522 ( .A(n10743), .B(n10799), .C(n5727), .Y(n2866) );
  OAI21X1 U1524 ( .A(n10743), .B(n10798), .C(n5993), .Y(n2867) );
  OAI21X1 U1526 ( .A(n10743), .B(n10797), .C(n5045), .Y(n2868) );
  OAI21X1 U1528 ( .A(n10744), .B(n10796), .C(n4936), .Y(n2869) );
  OAI21X1 U1530 ( .A(n10743), .B(n10795), .C(n5263), .Y(n2870) );
  OAI21X1 U1532 ( .A(n10743), .B(n10794), .C(n5155), .Y(n2871) );
  OAI21X1 U1534 ( .A(n10744), .B(n10793), .C(n5861), .Y(n2872) );
  OAI21X1 U1536 ( .A(n10743), .B(n10792), .C(n5372), .Y(n2873) );
  OAI21X1 U1538 ( .A(n10743), .B(n10791), .C(n6256), .Y(n2874) );
  OAI21X1 U1540 ( .A(n10743), .B(n10790), .C(n6124), .Y(n2875) );
  OAI21X1 U1542 ( .A(n10744), .B(n10789), .C(n5490), .Y(n2876) );
  OAI21X1 U1544 ( .A(n10744), .B(n10788), .C(n5154), .Y(n2877) );
  OAI21X1 U1546 ( .A(n10743), .B(n10787), .C(n5726), .Y(n2878) );
  OAI21X1 U1548 ( .A(n10744), .B(n10786), .C(n5044), .Y(n2879) );
  OAI21X1 U1550 ( .A(n10744), .B(n10785), .C(n5992), .Y(n2880) );
  OAI21X1 U1552 ( .A(n10743), .B(n10784), .C(n4618), .Y(n2881) );
  OAI21X1 U1554 ( .A(n10743), .B(n10783), .C(n5608), .Y(n2882) );
  OAI21X1 U1556 ( .A(n10743), .B(n10782), .C(n4512), .Y(n2883) );
  OAI21X1 U1558 ( .A(n10744), .B(n10781), .C(n4832), .Y(n2884) );
  OAI21X1 U1560 ( .A(n10744), .B(n10780), .C(n4725), .Y(n2885) );
  OAI21X1 U1562 ( .A(n10743), .B(n10779), .C(n4374), .Y(n2886) );
  OAI21X1 U1564 ( .A(n10744), .B(n10778), .C(n4373), .Y(n2887) );
  OAI21X1 U1566 ( .A(n10744), .B(n10777), .C(n4831), .Y(n2888) );
  OAI21X1 U1568 ( .A(n10743), .B(n10776), .C(n4372), .Y(n2889) );
  OAI21X1 U1570 ( .A(n10744), .B(n10775), .C(n4371), .Y(n2890) );
  OAI21X1 U1572 ( .A(n10744), .B(n10774), .C(n5262), .Y(n2891) );
  OAI21X1 U1574 ( .A(n10743), .B(n10773), .C(n4617), .Y(n2892) );
  OAI21X1 U1576 ( .A(n10744), .B(n10772), .C(n4511), .Y(n2893) );
  OAI21X1 U1578 ( .A(n10743), .B(n10771), .C(n5153), .Y(n2894) );
  OAI21X1 U1580 ( .A(n10743), .B(n10770), .C(n4370), .Y(n2895) );
  OAI21X1 U1582 ( .A(n10743), .B(n10769), .C(n4830), .Y(n2896) );
  OAI21X1 U1584 ( .A(n10744), .B(n10768), .C(n4369), .Y(n2897) );
  OAI21X1 U1586 ( .A(n10744), .B(n10767), .C(n4935), .Y(n2898) );
  OAI21X1 U1588 ( .A(n5772), .B(n6302), .C(reset_n), .Y(n827) );
  OAI21X1 U1589 ( .A(n10741), .B(n10830), .C(n5860), .Y(n2899) );
  OAI21X1 U1591 ( .A(n10741), .B(n10829), .C(n5859), .Y(n2900) );
  OAI21X1 U1593 ( .A(n10741), .B(n10828), .C(n5991), .Y(n2901) );
  OAI21X1 U1595 ( .A(n10741), .B(n10827), .C(n6123), .Y(n2902) );
  OAI21X1 U1597 ( .A(n10741), .B(n10826), .C(n6255), .Y(n2903) );
  OAI21X1 U1599 ( .A(n10741), .B(n10825), .C(n5371), .Y(n2904) );
  OAI21X1 U1601 ( .A(n10741), .B(n10824), .C(n5489), .Y(n2905) );
  OAI21X1 U1603 ( .A(n10741), .B(n10823), .C(n5607), .Y(n2906) );
  OAI21X1 U1605 ( .A(n10741), .B(n10822), .C(n5725), .Y(n2907) );
  OAI21X1 U1607 ( .A(n10741), .B(n10821), .C(n4934), .Y(n2908) );
  OAI21X1 U1609 ( .A(n10741), .B(n10820), .C(n5043), .Y(n2909) );
  OAI21X1 U1611 ( .A(n10741), .B(n10819), .C(n5152), .Y(n2910) );
  OAI21X1 U1613 ( .A(n10741), .B(n10818), .C(n5261), .Y(n2911) );
  OAI21X1 U1615 ( .A(n10741), .B(n10817), .C(n5858), .Y(n2912) );
  OAI21X1 U1617 ( .A(n10741), .B(n10816), .C(n5990), .Y(n2913) );
  OAI21X1 U1619 ( .A(n10741), .B(n10815), .C(n6122), .Y(n2914) );
  OAI21X1 U1621 ( .A(n10742), .B(n10814), .C(n6254), .Y(n2915) );
  OAI21X1 U1623 ( .A(n10742), .B(n10813), .C(n5370), .Y(n2916) );
  OAI21X1 U1625 ( .A(n10741), .B(n10812), .C(n5488), .Y(n2917) );
  OAI21X1 U1627 ( .A(n10742), .B(n10811), .C(n5606), .Y(n2918) );
  OAI21X1 U1629 ( .A(n10742), .B(n10810), .C(n5724), .Y(n2919) );
  OAI21X1 U1631 ( .A(n10742), .B(n10809), .C(n4933), .Y(n2920) );
  OAI21X1 U1633 ( .A(n10742), .B(n10808), .C(n5042), .Y(n2921) );
  OAI21X1 U1635 ( .A(n10741), .B(n10807), .C(n5151), .Y(n2922) );
  OAI21X1 U1637 ( .A(n10741), .B(n10806), .C(n4510), .Y(n2923) );
  OAI21X1 U1639 ( .A(n10741), .B(n10805), .C(n5723), .Y(n2924) );
  OAI21X1 U1641 ( .A(n10741), .B(n10804), .C(n5989), .Y(n2925) );
  OAI21X1 U1643 ( .A(n10741), .B(n10803), .C(n6121), .Y(n2926) );
  OAI21X1 U1645 ( .A(n10742), .B(n10802), .C(n6253), .Y(n2927) );
  OAI21X1 U1647 ( .A(n10741), .B(n10801), .C(n5369), .Y(n2928) );
  OAI21X1 U1649 ( .A(n10742), .B(n10800), .C(n5487), .Y(n2929) );
  OAI21X1 U1651 ( .A(n10741), .B(n10799), .C(n5605), .Y(n2930) );
  OAI21X1 U1653 ( .A(n10741), .B(n10798), .C(n5857), .Y(n2931) );
  OAI21X1 U1655 ( .A(n10741), .B(n10797), .C(n4932), .Y(n2932) );
  OAI21X1 U1657 ( .A(n10742), .B(n10796), .C(n5041), .Y(n2933) );
  OAI21X1 U1659 ( .A(n10741), .B(n10795), .C(n5150), .Y(n2934) );
  OAI21X1 U1661 ( .A(n10741), .B(n10794), .C(n5260), .Y(n2935) );
  OAI21X1 U1663 ( .A(n10742), .B(n10793), .C(n5988), .Y(n2936) );
  OAI21X1 U1665 ( .A(n10741), .B(n10792), .C(n5486), .Y(n2937) );
  OAI21X1 U1667 ( .A(n10741), .B(n10791), .C(n6120), .Y(n2938) );
  OAI21X1 U1669 ( .A(n10741), .B(n10790), .C(n6252), .Y(n2939) );
  OAI21X1 U1671 ( .A(n10742), .B(n10789), .C(n5368), .Y(n2940) );
  OAI21X1 U1673 ( .A(n10742), .B(n10788), .C(n5259), .Y(n2941) );
  OAI21X1 U1675 ( .A(n10741), .B(n10787), .C(n5604), .Y(n2942) );
  OAI21X1 U1677 ( .A(n10742), .B(n10786), .C(n4931), .Y(n2943) );
  OAI21X1 U1679 ( .A(n10742), .B(n10785), .C(n5856), .Y(n2944) );
  OAI21X1 U1681 ( .A(n10741), .B(n10784), .C(n4509), .Y(n2945) );
  OAI21X1 U1683 ( .A(n10741), .B(n10783), .C(n5722), .Y(n2946) );
  OAI21X1 U1685 ( .A(n10741), .B(n10782), .C(n4616), .Y(n2947) );
  OAI21X1 U1687 ( .A(n10742), .B(n10781), .C(n4724), .Y(n2948) );
  OAI21X1 U1689 ( .A(n10742), .B(n10780), .C(n4829), .Y(n2949) );
  OAI21X1 U1691 ( .A(n10741), .B(n10779), .C(n4368), .Y(n2950) );
  OAI21X1 U1693 ( .A(n10742), .B(n10778), .C(n4367), .Y(n2951) );
  OAI21X1 U1695 ( .A(n10742), .B(n10777), .C(n4723), .Y(n2952) );
  OAI21X1 U1697 ( .A(n10741), .B(n10776), .C(n4366), .Y(n2953) );
  OAI21X1 U1699 ( .A(n10742), .B(n10775), .C(n4365), .Y(n2954) );
  OAI21X1 U1701 ( .A(n10742), .B(n10774), .C(n5149), .Y(n2955) );
  OAI21X1 U1703 ( .A(n10741), .B(n10773), .C(n4508), .Y(n2956) );
  OAI21X1 U1705 ( .A(n10742), .B(n10772), .C(n4615), .Y(n2957) );
  OAI21X1 U1707 ( .A(n10741), .B(n10771), .C(n5258), .Y(n2958) );
  OAI21X1 U1709 ( .A(n10741), .B(n10770), .C(n4364), .Y(n2959) );
  OAI21X1 U1711 ( .A(n10741), .B(n10769), .C(n4722), .Y(n2960) );
  OAI21X1 U1713 ( .A(n10742), .B(n10768), .C(n4363), .Y(n2961) );
  OAI21X1 U1715 ( .A(n10742), .B(n10767), .C(n5040), .Y(n2962) );
  OAI21X1 U1717 ( .A(n5653), .B(n6302), .C(reset_n), .Y(n892) );
  OAI21X1 U1718 ( .A(n10739), .B(n10830), .C(n5721), .Y(n2963) );
  OAI21X1 U1720 ( .A(n10739), .B(n10829), .C(n5720), .Y(n2964) );
  OAI21X1 U1722 ( .A(n10739), .B(n10828), .C(n5603), .Y(n2965) );
  OAI21X1 U1724 ( .A(n10739), .B(n10827), .C(n5485), .Y(n2966) );
  OAI21X1 U1726 ( .A(n10739), .B(n10826), .C(n5367), .Y(n2967) );
  OAI21X1 U1728 ( .A(n10739), .B(n10825), .C(n6251), .Y(n2968) );
  OAI21X1 U1730 ( .A(n10739), .B(n10824), .C(n6119), .Y(n2969) );
  OAI21X1 U1732 ( .A(n10739), .B(n10823), .C(n5987), .Y(n2970) );
  OAI21X1 U1734 ( .A(n10739), .B(n10822), .C(n5855), .Y(n2971) );
  OAI21X1 U1736 ( .A(n10739), .B(n10821), .C(n4828), .Y(n2972) );
  OAI21X1 U1738 ( .A(n10739), .B(n10820), .C(n4721), .Y(n2973) );
  OAI21X1 U1740 ( .A(n10739), .B(n10819), .C(n4614), .Y(n2974) );
  OAI21X1 U1742 ( .A(n10739), .B(n10818), .C(n4507), .Y(n2975) );
  OAI21X1 U1744 ( .A(n10739), .B(n10817), .C(n5719), .Y(n2976) );
  OAI21X1 U1746 ( .A(n10739), .B(n10816), .C(n5602), .Y(n2977) );
  OAI21X1 U1748 ( .A(n10739), .B(n10815), .C(n5484), .Y(n2978) );
  OAI21X1 U1750 ( .A(n10740), .B(n10814), .C(n5366), .Y(n2979) );
  OAI21X1 U1752 ( .A(n10740), .B(n10813), .C(n6250), .Y(n2980) );
  OAI21X1 U1754 ( .A(n10739), .B(n10812), .C(n6118), .Y(n2981) );
  OAI21X1 U1756 ( .A(n10740), .B(n10811), .C(n5986), .Y(n2982) );
  OAI21X1 U1758 ( .A(n10740), .B(n10810), .C(n5854), .Y(n2983) );
  OAI21X1 U1760 ( .A(n10740), .B(n10809), .C(n4827), .Y(n2984) );
  OAI21X1 U1762 ( .A(n10740), .B(n10808), .C(n4720), .Y(n2985) );
  OAI21X1 U1764 ( .A(n10739), .B(n10807), .C(n4613), .Y(n2986) );
  OAI21X1 U1766 ( .A(n10739), .B(n10806), .C(n5257), .Y(n2987) );
  OAI21X1 U1768 ( .A(n10739), .B(n10805), .C(n5853), .Y(n2988) );
  OAI21X1 U1770 ( .A(n10739), .B(n10804), .C(n5601), .Y(n2989) );
  OAI21X1 U1772 ( .A(n10739), .B(n10803), .C(n5483), .Y(n2990) );
  OAI21X1 U1774 ( .A(n10740), .B(n10802), .C(n5365), .Y(n2991) );
  OAI21X1 U1776 ( .A(n10739), .B(n10801), .C(n6249), .Y(n2992) );
  OAI21X1 U1778 ( .A(n10740), .B(n10800), .C(n6117), .Y(n2993) );
  OAI21X1 U1780 ( .A(n10739), .B(n10799), .C(n5985), .Y(n2994) );
  OAI21X1 U1782 ( .A(n10739), .B(n10798), .C(n5718), .Y(n2995) );
  OAI21X1 U1784 ( .A(n10739), .B(n10797), .C(n4826), .Y(n2996) );
  OAI21X1 U1786 ( .A(n10740), .B(n10796), .C(n4719), .Y(n2997) );
  OAI21X1 U1788 ( .A(n10739), .B(n10795), .C(n4612), .Y(n2998) );
  OAI21X1 U1790 ( .A(n10739), .B(n10794), .C(n4506), .Y(n2999) );
  OAI21X1 U1792 ( .A(n10740), .B(n10793), .C(n5600), .Y(n3000) );
  OAI21X1 U1794 ( .A(n10739), .B(n10792), .C(n6116), .Y(n3001) );
  OAI21X1 U1796 ( .A(n10739), .B(n10791), .C(n5482), .Y(n3002) );
  OAI21X1 U1798 ( .A(n10739), .B(n10790), .C(n5364), .Y(n3003) );
  OAI21X1 U1800 ( .A(n10740), .B(n10789), .C(n6248), .Y(n3004) );
  OAI21X1 U1802 ( .A(n10740), .B(n10788), .C(n4505), .Y(n3005) );
  OAI21X1 U1804 ( .A(n10739), .B(n10787), .C(n5984), .Y(n3006) );
  OAI21X1 U1806 ( .A(n10740), .B(n10786), .C(n4825), .Y(n3007) );
  OAI21X1 U1808 ( .A(n10740), .B(n10785), .C(n5717), .Y(n3008) );
  OAI21X1 U1810 ( .A(n10739), .B(n10784), .C(n5256), .Y(n3009) );
  OAI21X1 U1812 ( .A(n10739), .B(n10783), .C(n5852), .Y(n3010) );
  OAI21X1 U1814 ( .A(n10739), .B(n10782), .C(n5148), .Y(n3011) );
  OAI21X1 U1816 ( .A(n10740), .B(n10781), .C(n5039), .Y(n3012) );
  OAI21X1 U1818 ( .A(n10740), .B(n10780), .C(n4930), .Y(n3013) );
  OAI21X1 U1820 ( .A(n10739), .B(n10779), .C(n4362), .Y(n3014) );
  OAI21X1 U1822 ( .A(n10740), .B(n10778), .C(n4361), .Y(n3015) );
  OAI21X1 U1824 ( .A(n10740), .B(n10777), .C(n5038), .Y(n3016) );
  OAI21X1 U1826 ( .A(n10739), .B(n10776), .C(n4360), .Y(n3017) );
  OAI21X1 U1828 ( .A(n10740), .B(n10775), .C(n4359), .Y(n3018) );
  OAI21X1 U1830 ( .A(n10740), .B(n10774), .C(n4611), .Y(n3019) );
  OAI21X1 U1832 ( .A(n10739), .B(n10773), .C(n5255), .Y(n3020) );
  OAI21X1 U1834 ( .A(n10740), .B(n10772), .C(n5147), .Y(n3021) );
  OAI21X1 U1836 ( .A(n10739), .B(n10771), .C(n4504), .Y(n3022) );
  OAI21X1 U1838 ( .A(n10739), .B(n10770), .C(n4358), .Y(n3023) );
  OAI21X1 U1840 ( .A(n10739), .B(n10769), .C(n5037), .Y(n3024) );
  OAI21X1 U1842 ( .A(n10740), .B(n10768), .C(n4357), .Y(n3025) );
  OAI21X1 U1844 ( .A(n10740), .B(n10767), .C(n4718), .Y(n3026) );
  OAI21X1 U1846 ( .A(n5771), .B(n6302), .C(reset_n), .Y(n957) );
  OAI21X1 U1847 ( .A(n10737), .B(n10830), .C(n5599), .Y(n3027) );
  OAI21X1 U1849 ( .A(n10737), .B(n10829), .C(n5598), .Y(n3028) );
  OAI21X1 U1851 ( .A(n10737), .B(n10828), .C(n5716), .Y(n3029) );
  OAI21X1 U1853 ( .A(n10737), .B(n10827), .C(n5363), .Y(n3030) );
  OAI21X1 U1855 ( .A(n10737), .B(n10826), .C(n5481), .Y(n3031) );
  OAI21X1 U1857 ( .A(n10737), .B(n10825), .C(n6115), .Y(n3032) );
  OAI21X1 U1859 ( .A(n10737), .B(n10824), .C(n6247), .Y(n3033) );
  OAI21X1 U1861 ( .A(n10737), .B(n10823), .C(n5851), .Y(n3034) );
  OAI21X1 U1863 ( .A(n10737), .B(n10822), .C(n5983), .Y(n3035) );
  OAI21X1 U1865 ( .A(n10737), .B(n10821), .C(n4717), .Y(n3036) );
  OAI21X1 U1867 ( .A(n10737), .B(n10820), .C(n4824), .Y(n3037) );
  OAI21X1 U1869 ( .A(n10737), .B(n10819), .C(n4503), .Y(n3038) );
  OAI21X1 U1871 ( .A(n10737), .B(n10818), .C(n4610), .Y(n3039) );
  OAI21X1 U1873 ( .A(n10737), .B(n10817), .C(n5597), .Y(n3040) );
  OAI21X1 U1875 ( .A(n10737), .B(n10816), .C(n5715), .Y(n3041) );
  OAI21X1 U1877 ( .A(n10737), .B(n10815), .C(n5362), .Y(n3042) );
  OAI21X1 U1879 ( .A(n10738), .B(n10814), .C(n5480), .Y(n3043) );
  OAI21X1 U1881 ( .A(n10738), .B(n10813), .C(n6114), .Y(n3044) );
  OAI21X1 U1883 ( .A(n10737), .B(n10812), .C(n6246), .Y(n3045) );
  OAI21X1 U1885 ( .A(n10738), .B(n10811), .C(n5850), .Y(n3046) );
  OAI21X1 U1887 ( .A(n10738), .B(n10810), .C(n5982), .Y(n3047) );
  OAI21X1 U1889 ( .A(n10738), .B(n10809), .C(n4716), .Y(n3048) );
  OAI21X1 U1891 ( .A(n10738), .B(n10808), .C(n4823), .Y(n3049) );
  OAI21X1 U1893 ( .A(n10737), .B(n10807), .C(n4502), .Y(n3050) );
  OAI21X1 U1895 ( .A(n10737), .B(n10806), .C(n5146), .Y(n3051) );
  OAI21X1 U1897 ( .A(n10737), .B(n10805), .C(n5981), .Y(n3052) );
  OAI21X1 U1899 ( .A(n10737), .B(n10804), .C(n5714), .Y(n3053) );
  OAI21X1 U1901 ( .A(n10737), .B(n10803), .C(n5361), .Y(n3054) );
  OAI21X1 U1903 ( .A(n10738), .B(n10802), .C(n5479), .Y(n3055) );
  OAI21X1 U1905 ( .A(n10737), .B(n10801), .C(n6113), .Y(n3056) );
  OAI21X1 U1907 ( .A(n10738), .B(n10800), .C(n6245), .Y(n3057) );
  OAI21X1 U1909 ( .A(n10737), .B(n10799), .C(n5849), .Y(n3058) );
  OAI21X1 U1911 ( .A(n10737), .B(n10798), .C(n5596), .Y(n3059) );
  OAI21X1 U1913 ( .A(n10737), .B(n10797), .C(n4715), .Y(n3060) );
  OAI21X1 U1915 ( .A(n10738), .B(n10796), .C(n4822), .Y(n3061) );
  OAI21X1 U1917 ( .A(n10737), .B(n10795), .C(n4501), .Y(n3062) );
  OAI21X1 U1919 ( .A(n10737), .B(n10794), .C(n4609), .Y(n3063) );
  OAI21X1 U1921 ( .A(n10738), .B(n10793), .C(n5713), .Y(n3064) );
  OAI21X1 U1923 ( .A(n10737), .B(n10792), .C(n6244), .Y(n3065) );
  OAI21X1 U1925 ( .A(n10737), .B(n10791), .C(n5360), .Y(n3066) );
  OAI21X1 U1927 ( .A(n10737), .B(n10790), .C(n5478), .Y(n3067) );
  OAI21X1 U1929 ( .A(n10738), .B(n10789), .C(n6112), .Y(n3068) );
  OAI21X1 U1931 ( .A(n10738), .B(n10788), .C(n4608), .Y(n3069) );
  OAI21X1 U1933 ( .A(n10737), .B(n10787), .C(n5848), .Y(n3070) );
  OAI21X1 U1935 ( .A(n10738), .B(n10786), .C(n4714), .Y(n3071) );
  OAI21X1 U1937 ( .A(n10738), .B(n10785), .C(n5595), .Y(n3072) );
  OAI21X1 U1939 ( .A(n10737), .B(n10784), .C(n5145), .Y(n3073) );
  OAI21X1 U1941 ( .A(n10737), .B(n10783), .C(n5980), .Y(n3074) );
  OAI21X1 U1943 ( .A(n10737), .B(n10782), .C(n5254), .Y(n3075) );
  OAI21X1 U1945 ( .A(n10738), .B(n10781), .C(n4929), .Y(n3076) );
  OAI21X1 U1947 ( .A(n10738), .B(n10780), .C(n5036), .Y(n3077) );
  OAI21X1 U1949 ( .A(n10737), .B(n10779), .C(n4356), .Y(n3078) );
  OAI21X1 U1951 ( .A(n10738), .B(n10778), .C(n4355), .Y(n3079) );
  OAI21X1 U1953 ( .A(n10738), .B(n10777), .C(n4928), .Y(n3080) );
  OAI21X1 U1955 ( .A(n10737), .B(n10776), .C(n4354), .Y(n3081) );
  OAI21X1 U1957 ( .A(n10738), .B(n10775), .C(n4353), .Y(n3082) );
  OAI21X1 U1959 ( .A(n10738), .B(n10774), .C(n4500), .Y(n3083) );
  OAI21X1 U1961 ( .A(n10737), .B(n10773), .C(n5144), .Y(n3084) );
  OAI21X1 U1963 ( .A(n10738), .B(n10772), .C(n5253), .Y(n3085) );
  OAI21X1 U1965 ( .A(n10737), .B(n10771), .C(n4607), .Y(n3086) );
  OAI21X1 U1967 ( .A(n10737), .B(n10770), .C(n4352), .Y(n3087) );
  OAI21X1 U1969 ( .A(n10737), .B(n10769), .C(n4927), .Y(n3088) );
  OAI21X1 U1971 ( .A(n10738), .B(n10768), .C(n4351), .Y(n3089) );
  OAI21X1 U1973 ( .A(n10738), .B(n10767), .C(n4821), .Y(n3090) );
  OAI21X1 U1975 ( .A(n5535), .B(n6302), .C(reset_n), .Y(n1022) );
  OAI21X1 U1976 ( .A(n10735), .B(n10830), .C(n5477), .Y(n3091) );
  OAI21X1 U1978 ( .A(n10735), .B(n10829), .C(n5476), .Y(n3092) );
  OAI21X1 U1980 ( .A(n10735), .B(n10828), .C(n5359), .Y(n3093) );
  OAI21X1 U1982 ( .A(n10735), .B(n10827), .C(n5712), .Y(n3094) );
  OAI21X1 U1984 ( .A(n10735), .B(n10826), .C(n5594), .Y(n3095) );
  OAI21X1 U1986 ( .A(n10735), .B(n10825), .C(n5979), .Y(n3096) );
  OAI21X1 U1988 ( .A(n10735), .B(n10824), .C(n5847), .Y(n3097) );
  OAI21X1 U1990 ( .A(n10735), .B(n10823), .C(n6243), .Y(n3098) );
  OAI21X1 U1992 ( .A(n10735), .B(n10822), .C(n6111), .Y(n3099) );
  OAI21X1 U1994 ( .A(n10735), .B(n10821), .C(n4606), .Y(n3100) );
  OAI21X1 U1996 ( .A(n10735), .B(n10820), .C(n4499), .Y(n3101) );
  OAI21X1 U1998 ( .A(n10735), .B(n10819), .C(n4820), .Y(n3102) );
  OAI21X1 U2000 ( .A(n10735), .B(n10818), .C(n4713), .Y(n3103) );
  OAI21X1 U2002 ( .A(n10735), .B(n10817), .C(n5475), .Y(n3104) );
  OAI21X1 U2004 ( .A(n10735), .B(n10816), .C(n5358), .Y(n3105) );
  OAI21X1 U2006 ( .A(n10735), .B(n10815), .C(n5711), .Y(n3106) );
  OAI21X1 U2008 ( .A(n10736), .B(n10814), .C(n5593), .Y(n3107) );
  OAI21X1 U2010 ( .A(n10736), .B(n10813), .C(n5978), .Y(n3108) );
  OAI21X1 U2012 ( .A(n10735), .B(n10812), .C(n5846), .Y(n3109) );
  OAI21X1 U2014 ( .A(n10736), .B(n10811), .C(n6242), .Y(n3110) );
  OAI21X1 U2016 ( .A(n10736), .B(n10810), .C(n6110), .Y(n3111) );
  OAI21X1 U2018 ( .A(n10736), .B(n10809), .C(n4605), .Y(n3112) );
  OAI21X1 U2020 ( .A(n10736), .B(n10808), .C(n4498), .Y(n3113) );
  OAI21X1 U2022 ( .A(n10735), .B(n10807), .C(n4819), .Y(n3114) );
  OAI21X1 U2024 ( .A(n10735), .B(n10806), .C(n5035), .Y(n3115) );
  OAI21X1 U2026 ( .A(n10735), .B(n10805), .C(n6109), .Y(n3116) );
  OAI21X1 U2028 ( .A(n10735), .B(n10804), .C(n5357), .Y(n3117) );
  OAI21X1 U2030 ( .A(n10735), .B(n10803), .C(n5710), .Y(n3118) );
  OAI21X1 U2032 ( .A(n10736), .B(n10802), .C(n5592), .Y(n3119) );
  OAI21X1 U2034 ( .A(n10735), .B(n10801), .C(n5977), .Y(n3120) );
  OAI21X1 U2036 ( .A(n10736), .B(n10800), .C(n5845), .Y(n3121) );
  OAI21X1 U2038 ( .A(n10735), .B(n10799), .C(n6241), .Y(n3122) );
  OAI21X1 U2040 ( .A(n10735), .B(n10798), .C(n5474), .Y(n3123) );
  OAI21X1 U2042 ( .A(n10735), .B(n10797), .C(n4604), .Y(n3124) );
  OAI21X1 U2044 ( .A(n10736), .B(n10796), .C(n4497), .Y(n3125) );
  OAI21X1 U2046 ( .A(n10735), .B(n10795), .C(n4818), .Y(n3126) );
  OAI21X1 U2048 ( .A(n10735), .B(n10794), .C(n4712), .Y(n3127) );
  OAI21X1 U2050 ( .A(n10736), .B(n10793), .C(n5356), .Y(n3128) );
  OAI21X1 U2052 ( .A(n10735), .B(n10792), .C(n5844), .Y(n3129) );
  OAI21X1 U2054 ( .A(n10735), .B(n10791), .C(n5709), .Y(n3130) );
  OAI21X1 U2056 ( .A(n10735), .B(n10790), .C(n5591), .Y(n3131) );
  OAI21X1 U2058 ( .A(n10736), .B(n10789), .C(n5976), .Y(n3132) );
  OAI21X1 U2060 ( .A(n10736), .B(n10788), .C(n4711), .Y(n3133) );
  OAI21X1 U2062 ( .A(n10735), .B(n10787), .C(n6240), .Y(n3134) );
  OAI21X1 U2064 ( .A(n10736), .B(n10786), .C(n4603), .Y(n3135) );
  OAI21X1 U2066 ( .A(n10736), .B(n10785), .C(n5473), .Y(n3136) );
  OAI21X1 U2068 ( .A(n10735), .B(n10784), .C(n5034), .Y(n3137) );
  OAI21X1 U2070 ( .A(n10735), .B(n10783), .C(n6108), .Y(n3138) );
  OAI21X1 U2072 ( .A(n10735), .B(n10782), .C(n4926), .Y(n3139) );
  OAI21X1 U2074 ( .A(n10736), .B(n10781), .C(n5252), .Y(n3140) );
  OAI21X1 U2076 ( .A(n10736), .B(n10780), .C(n5143), .Y(n3141) );
  OAI21X1 U2078 ( .A(n10735), .B(n10779), .C(n4350), .Y(n3142) );
  OAI21X1 U2080 ( .A(n10736), .B(n10778), .C(n4349), .Y(n3143) );
  OAI21X1 U2082 ( .A(n10736), .B(n10777), .C(n5251), .Y(n3144) );
  OAI21X1 U2084 ( .A(n10735), .B(n10776), .C(n4348), .Y(n3145) );
  OAI21X1 U2086 ( .A(n10736), .B(n10775), .C(n4347), .Y(n3146) );
  OAI21X1 U2088 ( .A(n10736), .B(n10774), .C(n4817), .Y(n3147) );
  OAI21X1 U2090 ( .A(n10735), .B(n10773), .C(n5033), .Y(n3148) );
  OAI21X1 U2092 ( .A(n10736), .B(n10772), .C(n4925), .Y(n3149) );
  OAI21X1 U2094 ( .A(n10735), .B(n10771), .C(n4710), .Y(n3150) );
  OAI21X1 U2096 ( .A(n10735), .B(n10770), .C(n4346), .Y(n3151) );
  OAI21X1 U2098 ( .A(n10735), .B(n10769), .C(n5250), .Y(n3152) );
  OAI21X1 U2100 ( .A(n10736), .B(n10768), .C(n4345), .Y(n3153) );
  OAI21X1 U2102 ( .A(n10736), .B(n10767), .C(n4496), .Y(n3154) );
  OAI21X1 U2104 ( .A(n5417), .B(n6302), .C(reset_n), .Y(n1087) );
  OAI21X1 U2105 ( .A(n10733), .B(n10830), .C(n5355), .Y(n3155) );
  OAI21X1 U2107 ( .A(n10733), .B(n10829), .C(n5354), .Y(n3156) );
  OAI21X1 U2109 ( .A(n10733), .B(n10828), .C(n5472), .Y(n3157) );
  OAI21X1 U2111 ( .A(n10733), .B(n10827), .C(n5590), .Y(n3158) );
  OAI21X1 U2113 ( .A(n10733), .B(n10826), .C(n5708), .Y(n3159) );
  OAI21X1 U2115 ( .A(n10733), .B(n10825), .C(n5843), .Y(n3160) );
  OAI21X1 U2117 ( .A(n10733), .B(n10824), .C(n5975), .Y(n3161) );
  OAI21X1 U2119 ( .A(n10733), .B(n10823), .C(n6107), .Y(n3162) );
  OAI21X1 U2121 ( .A(n10733), .B(n10822), .C(n6239), .Y(n3163) );
  OAI21X1 U2123 ( .A(n10733), .B(n10821), .C(n4495), .Y(n3164) );
  OAI21X1 U2125 ( .A(n10733), .B(n10820), .C(n4602), .Y(n3165) );
  OAI21X1 U2127 ( .A(n10733), .B(n10819), .C(n4709), .Y(n3166) );
  OAI21X1 U2129 ( .A(n10733), .B(n10818), .C(n4816), .Y(n3167) );
  OAI21X1 U2131 ( .A(n10733), .B(n10817), .C(n5353), .Y(n3168) );
  OAI21X1 U2133 ( .A(n10733), .B(n10816), .C(n5471), .Y(n3169) );
  OAI21X1 U2135 ( .A(n10734), .B(n10815), .C(n5589), .Y(n3170) );
  OAI21X1 U2137 ( .A(n10733), .B(n10814), .C(n5707), .Y(n3171) );
  OAI21X1 U2139 ( .A(n10734), .B(n10813), .C(n5842), .Y(n3172) );
  OAI21X1 U2141 ( .A(n10733), .B(n10812), .C(n5974), .Y(n3173) );
  OAI21X1 U2143 ( .A(n10734), .B(n10811), .C(n6106), .Y(n3174) );
  OAI21X1 U2145 ( .A(n10734), .B(n10810), .C(n6238), .Y(n3175) );
  OAI21X1 U2147 ( .A(n10734), .B(n10809), .C(n4494), .Y(n3176) );
  OAI21X1 U2149 ( .A(n10734), .B(n10808), .C(n4601), .Y(n3177) );
  OAI21X1 U2151 ( .A(n10733), .B(n10807), .C(n4708), .Y(n3178) );
  OAI21X1 U2153 ( .A(n10733), .B(n10806), .C(n4924), .Y(n3179) );
  OAI21X1 U2155 ( .A(n10733), .B(n10805), .C(n6237), .Y(n3180) );
  OAI21X1 U2157 ( .A(n10733), .B(n10804), .C(n5470), .Y(n3181) );
  OAI21X1 U2159 ( .A(n10733), .B(n10803), .C(n5588), .Y(n3182) );
  OAI21X1 U2161 ( .A(n10734), .B(n10802), .C(n5706), .Y(n3183) );
  OAI21X1 U2163 ( .A(n10734), .B(n10801), .C(n5841), .Y(n3184) );
  OAI21X1 U2165 ( .A(n10734), .B(n10800), .C(n5973), .Y(n3185) );
  OAI21X1 U2167 ( .A(n10733), .B(n10799), .C(n6105), .Y(n3186) );
  OAI21X1 U2169 ( .A(n10733), .B(n10798), .C(n5352), .Y(n3187) );
  OAI21X1 U2171 ( .A(n10733), .B(n10797), .C(n4493), .Y(n3188) );
  OAI21X1 U2173 ( .A(n10733), .B(n10796), .C(n4600), .Y(n3189) );
  OAI21X1 U2175 ( .A(n10734), .B(n10795), .C(n4707), .Y(n3190) );
  OAI21X1 U2177 ( .A(n10733), .B(n10794), .C(n4815), .Y(n3191) );
  OAI21X1 U2179 ( .A(n10733), .B(n10793), .C(n5469), .Y(n3192) );
  OAI21X1 U2181 ( .A(n10733), .B(n10792), .C(n5972), .Y(n3193) );
  OAI21X1 U2183 ( .A(n10733), .B(n10791), .C(n5587), .Y(n3194) );
  OAI21X1 U2185 ( .A(n10733), .B(n10790), .C(n5705), .Y(n3195) );
  OAI21X1 U2187 ( .A(n10734), .B(n10789), .C(n5840), .Y(n3196) );
  OAI21X1 U2189 ( .A(n10734), .B(n10788), .C(n4814), .Y(n3197) );
  OAI21X1 U2191 ( .A(n10733), .B(n10787), .C(n6104), .Y(n3198) );
  OAI21X1 U2193 ( .A(n10734), .B(n10786), .C(n4492), .Y(n3199) );
  OAI21X1 U2195 ( .A(n10734), .B(n10785), .C(n5351), .Y(n3200) );
  OAI21X1 U2197 ( .A(n10733), .B(n10784), .C(n4923), .Y(n3201) );
  OAI21X1 U2199 ( .A(n10734), .B(n10783), .C(n6236), .Y(n3202) );
  OAI21X1 U2201 ( .A(n10733), .B(n10782), .C(n5032), .Y(n3203) );
  OAI21X1 U2203 ( .A(n10734), .B(n10781), .C(n5142), .Y(n3204) );
  OAI21X1 U2205 ( .A(n10734), .B(n10780), .C(n5249), .Y(n3205) );
  OAI21X1 U2207 ( .A(n10734), .B(n10779), .C(n4344), .Y(n3206) );
  OAI21X1 U2209 ( .A(n10733), .B(n10778), .C(n4343), .Y(n3207) );
  OAI21X1 U2211 ( .A(n10733), .B(n10777), .C(n5141), .Y(n3208) );
  OAI21X1 U2213 ( .A(n10733), .B(n10776), .C(n4342), .Y(n3209) );
  OAI21X1 U2215 ( .A(n10734), .B(n10775), .C(n4341), .Y(n3210) );
  OAI21X1 U2217 ( .A(n10734), .B(n10774), .C(n4706), .Y(n3211) );
  OAI21X1 U2219 ( .A(n10733), .B(n10773), .C(n4922), .Y(n3212) );
  OAI21X1 U2221 ( .A(n10734), .B(n10772), .C(n5031), .Y(n3213) );
  OAI21X1 U2223 ( .A(n10733), .B(n10771), .C(n4813), .Y(n3214) );
  OAI21X1 U2225 ( .A(n10733), .B(n10770), .C(n4340), .Y(n3215) );
  OAI21X1 U2227 ( .A(n10733), .B(n10769), .C(n5140), .Y(n3216) );
  OAI21X1 U2229 ( .A(n10734), .B(n10768), .C(n4339), .Y(n3217) );
  OAI21X1 U2231 ( .A(n10734), .B(n10767), .C(n4599), .Y(n3218) );
  OAI21X1 U2233 ( .A(n5299), .B(n6302), .C(reset_n), .Y(n1152) );
  NAND3X1 U2234 ( .A(n10765), .B(n10832), .C(waddr[4]), .Y(n697) );
  OAI21X1 U2235 ( .A(n10731), .B(n10830), .C(n5248), .Y(n3219) );
  OAI21X1 U2237 ( .A(n10731), .B(n10829), .C(n5247), .Y(n3220) );
  OAI21X1 U2239 ( .A(n10731), .B(n10828), .C(n5139), .Y(n3221) );
  OAI21X1 U2241 ( .A(n10731), .B(n10827), .C(n5030), .Y(n3222) );
  OAI21X1 U2243 ( .A(n10731), .B(n10826), .C(n4921), .Y(n3223) );
  OAI21X1 U2245 ( .A(n10731), .B(n10825), .C(n4812), .Y(n3224) );
  OAI21X1 U2247 ( .A(n10731), .B(n10824), .C(n4705), .Y(n3225) );
  OAI21X1 U2249 ( .A(n10731), .B(n10823), .C(n4598), .Y(n3226) );
  OAI21X1 U2251 ( .A(n10731), .B(n10822), .C(n4491), .Y(n3227) );
  OAI21X1 U2253 ( .A(n10731), .B(n10821), .C(n6235), .Y(n3228) );
  OAI21X1 U2255 ( .A(n10731), .B(n10820), .C(n6103), .Y(n3229) );
  OAI21X1 U2257 ( .A(n10731), .B(n10819), .C(n5971), .Y(n3230) );
  OAI21X1 U2259 ( .A(n10731), .B(n10818), .C(n5839), .Y(n3231) );
  OAI21X1 U2261 ( .A(n10731), .B(n10817), .C(n5246), .Y(n3232) );
  OAI21X1 U2263 ( .A(n10731), .B(n10816), .C(n5138), .Y(n3233) );
  OAI21X1 U2265 ( .A(n10732), .B(n10815), .C(n5029), .Y(n3234) );
  OAI21X1 U2267 ( .A(n10731), .B(n10814), .C(n4920), .Y(n3235) );
  OAI21X1 U2269 ( .A(n10732), .B(n10813), .C(n4811), .Y(n3236) );
  OAI21X1 U2271 ( .A(n10731), .B(n10812), .C(n4704), .Y(n3237) );
  OAI21X1 U2273 ( .A(n10732), .B(n10811), .C(n4597), .Y(n3238) );
  OAI21X1 U2275 ( .A(n10732), .B(n10810), .C(n4490), .Y(n3239) );
  OAI21X1 U2277 ( .A(n10732), .B(n10809), .C(n6234), .Y(n3240) );
  OAI21X1 U2279 ( .A(n10732), .B(n10808), .C(n6102), .Y(n3241) );
  OAI21X1 U2281 ( .A(n10731), .B(n10807), .C(n5970), .Y(n3242) );
  OAI21X1 U2283 ( .A(n10731), .B(n10806), .C(n5704), .Y(n3243) );
  OAI21X1 U2285 ( .A(n10731), .B(n10805), .C(n4489), .Y(n3244) );
  OAI21X1 U2287 ( .A(n10731), .B(n10804), .C(n5137), .Y(n3245) );
  OAI21X1 U2289 ( .A(n10731), .B(n10803), .C(n5028), .Y(n3246) );
  OAI21X1 U2291 ( .A(n10732), .B(n10802), .C(n4919), .Y(n3247) );
  OAI21X1 U2293 ( .A(n10732), .B(n10801), .C(n4810), .Y(n3248) );
  OAI21X1 U2295 ( .A(n10732), .B(n10800), .C(n4703), .Y(n3249) );
  OAI21X1 U2297 ( .A(n10731), .B(n10799), .C(n4596), .Y(n3250) );
  OAI21X1 U2299 ( .A(n10731), .B(n10798), .C(n5245), .Y(n3251) );
  OAI21X1 U2301 ( .A(n10731), .B(n10797), .C(n6233), .Y(n3252) );
  OAI21X1 U2303 ( .A(n10731), .B(n10796), .C(n6101), .Y(n3253) );
  OAI21X1 U2305 ( .A(n10732), .B(n10795), .C(n5969), .Y(n3254) );
  OAI21X1 U2307 ( .A(n10731), .B(n10794), .C(n5838), .Y(n3255) );
  OAI21X1 U2309 ( .A(n10731), .B(n10793), .C(n5136), .Y(n3256) );
  OAI21X1 U2311 ( .A(n10731), .B(n10792), .C(n4702), .Y(n3257) );
  OAI21X1 U2313 ( .A(n10731), .B(n10791), .C(n5027), .Y(n3258) );
  OAI21X1 U2315 ( .A(n10731), .B(n10790), .C(n4918), .Y(n3259) );
  OAI21X1 U2317 ( .A(n10732), .B(n10789), .C(n4809), .Y(n3260) );
  OAI21X1 U2319 ( .A(n10732), .B(n10788), .C(n5837), .Y(n3261) );
  OAI21X1 U2321 ( .A(n10731), .B(n10787), .C(n4595), .Y(n3262) );
  OAI21X1 U2323 ( .A(n10732), .B(n10786), .C(n6232), .Y(n3263) );
  OAI21X1 U2325 ( .A(n10732), .B(n10785), .C(n5244), .Y(n3264) );
  OAI21X1 U2327 ( .A(n10731), .B(n10784), .C(n5703), .Y(n3265) );
  OAI21X1 U2329 ( .A(n10732), .B(n10783), .C(n4488), .Y(n3266) );
  OAI21X1 U2331 ( .A(n10731), .B(n10782), .C(n5586), .Y(n3267) );
  OAI21X1 U2333 ( .A(n10732), .B(n10781), .C(n5468), .Y(n3268) );
  OAI21X1 U2335 ( .A(n10732), .B(n10780), .C(n5350), .Y(n3269) );
  OAI21X1 U2337 ( .A(n10732), .B(n10779), .C(n4338), .Y(n3270) );
  OAI21X1 U2339 ( .A(n10731), .B(n10778), .C(n4337), .Y(n3271) );
  OAI21X1 U2341 ( .A(n10731), .B(n10777), .C(n5467), .Y(n3272) );
  OAI21X1 U2343 ( .A(n10731), .B(n10776), .C(n4336), .Y(n3273) );
  OAI21X1 U2345 ( .A(n10732), .B(n10775), .C(n4335), .Y(n3274) );
  OAI21X1 U2347 ( .A(n10732), .B(n10774), .C(n5968), .Y(n3275) );
  OAI21X1 U2349 ( .A(n10731), .B(n10773), .C(n5702), .Y(n3276) );
  OAI21X1 U2351 ( .A(n10732), .B(n10772), .C(n5585), .Y(n3277) );
  OAI21X1 U2353 ( .A(n10731), .B(n10771), .C(n5836), .Y(n3278) );
  OAI21X1 U2355 ( .A(n10731), .B(n10770), .C(n4334), .Y(n3279) );
  OAI21X1 U2357 ( .A(n10731), .B(n10769), .C(n5466), .Y(n3280) );
  OAI21X1 U2359 ( .A(n10732), .B(n10768), .C(n4333), .Y(n3281) );
  OAI21X1 U2361 ( .A(n10732), .B(n10767), .C(n6100), .Y(n3282) );
  OAI21X1 U2363 ( .A(n5774), .B(n6170), .C(reset_n), .Y(n1217) );
  OAI21X1 U2364 ( .A(n10729), .B(n10830), .C(n5135), .Y(n3283) );
  OAI21X1 U2366 ( .A(n10729), .B(n10829), .C(n5134), .Y(n3284) );
  OAI21X1 U2368 ( .A(n10729), .B(n10828), .C(n5243), .Y(n3285) );
  OAI21X1 U2370 ( .A(n10729), .B(n10827), .C(n4917), .Y(n3286) );
  OAI21X1 U2372 ( .A(n10729), .B(n10826), .C(n5026), .Y(n3287) );
  OAI21X1 U2374 ( .A(n10729), .B(n10825), .C(n4701), .Y(n3288) );
  OAI21X1 U2376 ( .A(n10729), .B(n10824), .C(n4808), .Y(n3289) );
  OAI21X1 U2378 ( .A(n10729), .B(n10823), .C(n4487), .Y(n3290) );
  OAI21X1 U2380 ( .A(n10729), .B(n10822), .C(n4594), .Y(n3291) );
  OAI21X1 U2382 ( .A(n10729), .B(n10821), .C(n6099), .Y(n3292) );
  OAI21X1 U2384 ( .A(n10729), .B(n10820), .C(n6231), .Y(n3293) );
  OAI21X1 U2386 ( .A(n10729), .B(n10819), .C(n5835), .Y(n3294) );
  OAI21X1 U2388 ( .A(n10729), .B(n10818), .C(n5967), .Y(n3295) );
  OAI21X1 U2390 ( .A(n10729), .B(n10817), .C(n5133), .Y(n3296) );
  OAI21X1 U2392 ( .A(n10729), .B(n10816), .C(n5242), .Y(n3297) );
  OAI21X1 U2394 ( .A(n10729), .B(n10815), .C(n4916), .Y(n3298) );
  OAI21X1 U2396 ( .A(n10730), .B(n10814), .C(n5025), .Y(n3299) );
  OAI21X1 U2398 ( .A(n10730), .B(n10813), .C(n4700), .Y(n3300) );
  OAI21X1 U2400 ( .A(n10729), .B(n10812), .C(n4807), .Y(n3301) );
  OAI21X1 U2402 ( .A(n10730), .B(n10811), .C(n4486), .Y(n3302) );
  OAI21X1 U2404 ( .A(n10730), .B(n10810), .C(n4593), .Y(n3303) );
  OAI21X1 U2406 ( .A(n10730), .B(n10809), .C(n6098), .Y(n3304) );
  OAI21X1 U2408 ( .A(n10730), .B(n10808), .C(n6230), .Y(n3305) );
  OAI21X1 U2410 ( .A(n10729), .B(n10807), .C(n5834), .Y(n3306) );
  OAI21X1 U2412 ( .A(n10729), .B(n10806), .C(n5584), .Y(n3307) );
  OAI21X1 U2414 ( .A(n10729), .B(n10805), .C(n4592), .Y(n3308) );
  OAI21X1 U2416 ( .A(n10729), .B(n10804), .C(n5241), .Y(n3309) );
  OAI21X1 U2418 ( .A(n10729), .B(n10803), .C(n4915), .Y(n3310) );
  OAI21X1 U2420 ( .A(n10730), .B(n10802), .C(n5024), .Y(n3311) );
  OAI21X1 U2422 ( .A(n10729), .B(n10801), .C(n4699), .Y(n3312) );
  OAI21X1 U2424 ( .A(n10730), .B(n10800), .C(n4806), .Y(n3313) );
  OAI21X1 U2426 ( .A(n10729), .B(n10799), .C(n4485), .Y(n3314) );
  OAI21X1 U2428 ( .A(n10729), .B(n10798), .C(n5132), .Y(n3315) );
  OAI21X1 U2430 ( .A(n10729), .B(n10797), .C(n6097), .Y(n3316) );
  OAI21X1 U2432 ( .A(n10730), .B(n10796), .C(n6229), .Y(n3317) );
  OAI21X1 U2434 ( .A(n10729), .B(n10795), .C(n5833), .Y(n3318) );
  OAI21X1 U2436 ( .A(n10729), .B(n10794), .C(n5966), .Y(n3319) );
  OAI21X1 U2438 ( .A(n10730), .B(n10793), .C(n5240), .Y(n3320) );
  OAI21X1 U2440 ( .A(n10729), .B(n10792), .C(n4805), .Y(n3321) );
  OAI21X1 U2442 ( .A(n10729), .B(n10791), .C(n4914), .Y(n3322) );
  OAI21X1 U2444 ( .A(n10729), .B(n10790), .C(n5023), .Y(n3323) );
  OAI21X1 U2446 ( .A(n10730), .B(n10789), .C(n4698), .Y(n3324) );
  OAI21X1 U2448 ( .A(n10730), .B(n10788), .C(n5965), .Y(n3325) );
  OAI21X1 U2450 ( .A(n10729), .B(n10787), .C(n4484), .Y(n3326) );
  OAI21X1 U2452 ( .A(n10730), .B(n10786), .C(n6096), .Y(n3327) );
  OAI21X1 U2454 ( .A(n10730), .B(n10785), .C(n5131), .Y(n3328) );
  OAI21X1 U2456 ( .A(n10729), .B(n10784), .C(n5583), .Y(n3329) );
  OAI21X1 U2458 ( .A(n10729), .B(n10783), .C(n4591), .Y(n3330) );
  OAI21X1 U2460 ( .A(n10729), .B(n10782), .C(n5701), .Y(n3331) );
  OAI21X1 U2462 ( .A(n10730), .B(n10781), .C(n5349), .Y(n3332) );
  OAI21X1 U2464 ( .A(n10730), .B(n10780), .C(n5465), .Y(n3333) );
  OAI21X1 U2466 ( .A(n10729), .B(n10779), .C(n4332), .Y(n3334) );
  OAI21X1 U2468 ( .A(n10730), .B(n10778), .C(n4331), .Y(n3335) );
  OAI21X1 U2470 ( .A(n10730), .B(n10777), .C(n5348), .Y(n3336) );
  OAI21X1 U2472 ( .A(n10729), .B(n10776), .C(n4330), .Y(n3337) );
  OAI21X1 U2474 ( .A(n10730), .B(n10775), .C(n4329), .Y(n3338) );
  OAI21X1 U2476 ( .A(n10730), .B(n10774), .C(n5832), .Y(n3339) );
  OAI21X1 U2478 ( .A(n10729), .B(n10773), .C(n5582), .Y(n3340) );
  OAI21X1 U2480 ( .A(n10730), .B(n10772), .C(n5700), .Y(n3341) );
  OAI21X1 U2482 ( .A(n10729), .B(n10771), .C(n5964), .Y(n3342) );
  OAI21X1 U2484 ( .A(n10729), .B(n10770), .C(n4328), .Y(n3343) );
  OAI21X1 U2486 ( .A(n10729), .B(n10769), .C(n5347), .Y(n3344) );
  OAI21X1 U2488 ( .A(n10730), .B(n10768), .C(n4327), .Y(n3345) );
  OAI21X1 U2490 ( .A(n10730), .B(n10767), .C(n6228), .Y(n3346) );
  OAI21X1 U2492 ( .A(n5773), .B(n6170), .C(reset_n), .Y(n1283) );
  OAI21X1 U2493 ( .A(n10727), .B(n10830), .C(n5022), .Y(n3347) );
  OAI21X1 U2495 ( .A(n10727), .B(n10829), .C(n5021), .Y(n3348) );
  OAI21X1 U2497 ( .A(n10727), .B(n10828), .C(n4913), .Y(n3349) );
  OAI21X1 U2499 ( .A(n10727), .B(n10827), .C(n5239), .Y(n3350) );
  OAI21X1 U2501 ( .A(n10727), .B(n10826), .C(n5130), .Y(n3351) );
  OAI21X1 U2503 ( .A(n10727), .B(n10825), .C(n4590), .Y(n3352) );
  OAI21X1 U2505 ( .A(n10727), .B(n10824), .C(n4483), .Y(n3353) );
  OAI21X1 U2507 ( .A(n10727), .B(n10823), .C(n4804), .Y(n3354) );
  OAI21X1 U2509 ( .A(n10727), .B(n10822), .C(n4697), .Y(n3355) );
  OAI21X1 U2511 ( .A(n10727), .B(n10821), .C(n5963), .Y(n3356) );
  OAI21X1 U2513 ( .A(n10727), .B(n10820), .C(n5831), .Y(n3357) );
  OAI21X1 U2515 ( .A(n10727), .B(n10819), .C(n6227), .Y(n3358) );
  OAI21X1 U2517 ( .A(n10727), .B(n10818), .C(n6095), .Y(n3359) );
  OAI21X1 U2519 ( .A(n10727), .B(n10817), .C(n5020), .Y(n3360) );
  OAI21X1 U2521 ( .A(n10727), .B(n10816), .C(n4912), .Y(n3361) );
  OAI21X1 U2523 ( .A(n10728), .B(n10815), .C(n5238), .Y(n3362) );
  OAI21X1 U2525 ( .A(n10727), .B(n10814), .C(n5129), .Y(n3363) );
  OAI21X1 U2527 ( .A(n10728), .B(n10813), .C(n4589), .Y(n3364) );
  OAI21X1 U2529 ( .A(n10727), .B(n10812), .C(n4482), .Y(n3365) );
  OAI21X1 U2531 ( .A(n10728), .B(n10811), .C(n4803), .Y(n3366) );
  OAI21X1 U2533 ( .A(n10728), .B(n10810), .C(n4696), .Y(n3367) );
  OAI21X1 U2535 ( .A(n10728), .B(n10809), .C(n5962), .Y(n3368) );
  OAI21X1 U2537 ( .A(n10728), .B(n10808), .C(n5830), .Y(n3369) );
  OAI21X1 U2539 ( .A(n10727), .B(n10807), .C(n6226), .Y(n3370) );
  OAI21X1 U2541 ( .A(n10727), .B(n10806), .C(n5464), .Y(n3371) );
  OAI21X1 U2543 ( .A(n10727), .B(n10805), .C(n4695), .Y(n3372) );
  OAI21X1 U2545 ( .A(n10727), .B(n10804), .C(n4911), .Y(n3373) );
  OAI21X1 U2547 ( .A(n10727), .B(n10803), .C(n5237), .Y(n3374) );
  OAI21X1 U2549 ( .A(n10728), .B(n10802), .C(n5128), .Y(n3375) );
  OAI21X1 U2551 ( .A(n10728), .B(n10801), .C(n4588), .Y(n3376) );
  OAI21X1 U2553 ( .A(n10728), .B(n10800), .C(n4481), .Y(n3377) );
  OAI21X1 U2555 ( .A(n10727), .B(n10799), .C(n4802), .Y(n3378) );
  OAI21X1 U2557 ( .A(n10727), .B(n10798), .C(n5019), .Y(n3379) );
  OAI21X1 U2559 ( .A(n10727), .B(n10797), .C(n5961), .Y(n3380) );
  OAI21X1 U2561 ( .A(n10727), .B(n10796), .C(n5829), .Y(n3381) );
  OAI21X1 U2563 ( .A(n10728), .B(n10795), .C(n6225), .Y(n3382) );
  OAI21X1 U2565 ( .A(n10727), .B(n10794), .C(n6094), .Y(n3383) );
  OAI21X1 U2567 ( .A(n10727), .B(n10793), .C(n4910), .Y(n3384) );
  OAI21X1 U2569 ( .A(n10727), .B(n10792), .C(n4480), .Y(n3385) );
  OAI21X1 U2571 ( .A(n10727), .B(n10791), .C(n5236), .Y(n3386) );
  OAI21X1 U2573 ( .A(n10727), .B(n10790), .C(n5127), .Y(n3387) );
  OAI21X1 U2575 ( .A(n10728), .B(n10789), .C(n4587), .Y(n3388) );
  OAI21X1 U2577 ( .A(n10728), .B(n10788), .C(n6093), .Y(n3389) );
  OAI21X1 U2579 ( .A(n10727), .B(n10787), .C(n4801), .Y(n3390) );
  OAI21X1 U2581 ( .A(n10728), .B(n10786), .C(n5960), .Y(n3391) );
  OAI21X1 U2583 ( .A(n10728), .B(n10785), .C(n5018), .Y(n3392) );
  OAI21X1 U2585 ( .A(n10727), .B(n10784), .C(n5463), .Y(n3393) );
  OAI21X1 U2587 ( .A(n10728), .B(n10783), .C(n4694), .Y(n3394) );
  OAI21X1 U2589 ( .A(n10727), .B(n10782), .C(n5346), .Y(n3395) );
  OAI21X1 U2591 ( .A(n10728), .B(n10781), .C(n5699), .Y(n3396) );
  OAI21X1 U2593 ( .A(n10728), .B(n10780), .C(n5581), .Y(n3397) );
  OAI21X1 U2595 ( .A(n10728), .B(n10779), .C(n4326), .Y(n3398) );
  OAI21X1 U2597 ( .A(n10727), .B(n10778), .C(n4325), .Y(n3399) );
  OAI21X1 U2599 ( .A(n10727), .B(n10777), .C(n5698), .Y(n3400) );
  OAI21X1 U2601 ( .A(n10727), .B(n10776), .C(n4324), .Y(n3401) );
  OAI21X1 U2603 ( .A(n10728), .B(n10775), .C(n4323), .Y(n3402) );
  OAI21X1 U2605 ( .A(n10728), .B(n10774), .C(n6224), .Y(n3403) );
  OAI21X1 U2607 ( .A(n10727), .B(n10773), .C(n5462), .Y(n3404) );
  OAI21X1 U2609 ( .A(n10728), .B(n10772), .C(n5345), .Y(n3405) );
  OAI21X1 U2611 ( .A(n10727), .B(n10771), .C(n6092), .Y(n3406) );
  OAI21X1 U2613 ( .A(n10727), .B(n10770), .C(n4322), .Y(n3407) );
  OAI21X1 U2615 ( .A(n10727), .B(n10769), .C(n5697), .Y(n3408) );
  OAI21X1 U2617 ( .A(n10728), .B(n10768), .C(n4321), .Y(n3409) );
  OAI21X1 U2619 ( .A(n10728), .B(n10767), .C(n5828), .Y(n3410) );
  OAI21X1 U2621 ( .A(n5772), .B(n6170), .C(reset_n), .Y(n1348) );
  OAI21X1 U2622 ( .A(n10725), .B(n10830), .C(n4909), .Y(n3411) );
  OAI21X1 U2624 ( .A(n10725), .B(n10829), .C(n4908), .Y(n3412) );
  OAI21X1 U2626 ( .A(n10725), .B(n10828), .C(n5017), .Y(n3413) );
  OAI21X1 U2628 ( .A(n10725), .B(n10827), .C(n5126), .Y(n3414) );
  OAI21X1 U2630 ( .A(n10725), .B(n10826), .C(n5235), .Y(n3415) );
  OAI21X1 U2632 ( .A(n10725), .B(n10825), .C(n4479), .Y(n3416) );
  OAI21X1 U2634 ( .A(n10725), .B(n10824), .C(n4586), .Y(n3417) );
  OAI21X1 U2636 ( .A(n10725), .B(n10823), .C(n4693), .Y(n3418) );
  OAI21X1 U2638 ( .A(n10725), .B(n10822), .C(n4800), .Y(n3419) );
  OAI21X1 U2640 ( .A(n10725), .B(n10821), .C(n5827), .Y(n3420) );
  OAI21X1 U2642 ( .A(n10725), .B(n10820), .C(n5959), .Y(n3421) );
  OAI21X1 U2644 ( .A(n10725), .B(n10819), .C(n6091), .Y(n3422) );
  OAI21X1 U2646 ( .A(n10725), .B(n10818), .C(n6223), .Y(n3423) );
  OAI21X1 U2648 ( .A(n10725), .B(n10817), .C(n4907), .Y(n3424) );
  OAI21X1 U2650 ( .A(n10725), .B(n10816), .C(n5016), .Y(n3425) );
  OAI21X1 U2652 ( .A(n10726), .B(n10815), .C(n5125), .Y(n3426) );
  OAI21X1 U2654 ( .A(n10725), .B(n10814), .C(n5234), .Y(n3427) );
  OAI21X1 U2656 ( .A(n10726), .B(n10813), .C(n4478), .Y(n3428) );
  OAI21X1 U2658 ( .A(n10725), .B(n10812), .C(n4585), .Y(n3429) );
  OAI21X1 U2660 ( .A(n10726), .B(n10811), .C(n4692), .Y(n3430) );
  OAI21X1 U2662 ( .A(n10726), .B(n10810), .C(n4799), .Y(n3431) );
  OAI21X1 U2664 ( .A(n10726), .B(n10809), .C(n5826), .Y(n3432) );
  OAI21X1 U2666 ( .A(n10726), .B(n10808), .C(n5958), .Y(n3433) );
  OAI21X1 U2668 ( .A(n10725), .B(n10807), .C(n6090), .Y(n3434) );
  OAI21X1 U2670 ( .A(n10725), .B(n10806), .C(n5344), .Y(n3435) );
  OAI21X1 U2672 ( .A(n10725), .B(n10805), .C(n4798), .Y(n3436) );
  OAI21X1 U2674 ( .A(n10725), .B(n10804), .C(n5015), .Y(n3437) );
  OAI21X1 U2676 ( .A(n10725), .B(n10803), .C(n5124), .Y(n3438) );
  OAI21X1 U2678 ( .A(n10726), .B(n10802), .C(n5233), .Y(n3439) );
  OAI21X1 U2680 ( .A(n10726), .B(n10801), .C(n4477), .Y(n3440) );
  OAI21X1 U2682 ( .A(n10726), .B(n10800), .C(n4584), .Y(n3441) );
  OAI21X1 U2684 ( .A(n10725), .B(n10799), .C(n4691), .Y(n3442) );
  OAI21X1 U2686 ( .A(n10725), .B(n10798), .C(n4906), .Y(n3443) );
  OAI21X1 U2688 ( .A(n10725), .B(n10797), .C(n5825), .Y(n3444) );
  OAI21X1 U2690 ( .A(n10725), .B(n10796), .C(n5957), .Y(n3445) );
  OAI21X1 U2692 ( .A(n10726), .B(n10795), .C(n6089), .Y(n3446) );
  OAI21X1 U2694 ( .A(n10725), .B(n10794), .C(n6222), .Y(n3447) );
  OAI21X1 U2696 ( .A(n10725), .B(n10793), .C(n5014), .Y(n3448) );
  OAI21X1 U2698 ( .A(n10725), .B(n10792), .C(n4583), .Y(n3449) );
  OAI21X1 U2700 ( .A(n10725), .B(n10791), .C(n5123), .Y(n3450) );
  OAI21X1 U2702 ( .A(n10725), .B(n10790), .C(n5232), .Y(n3451) );
  OAI21X1 U2704 ( .A(n10726), .B(n10789), .C(n4476), .Y(n3452) );
  OAI21X1 U2706 ( .A(n10726), .B(n10788), .C(n6221), .Y(n3453) );
  OAI21X1 U2708 ( .A(n10725), .B(n10787), .C(n4690), .Y(n3454) );
  OAI21X1 U2710 ( .A(n10726), .B(n10786), .C(n5824), .Y(n3455) );
  OAI21X1 U2712 ( .A(n10726), .B(n10785), .C(n4905), .Y(n3456) );
  OAI21X1 U2714 ( .A(n10725), .B(n10784), .C(n5343), .Y(n3457) );
  OAI21X1 U2716 ( .A(n10726), .B(n10783), .C(n4797), .Y(n3458) );
  OAI21X1 U2718 ( .A(n10725), .B(n10782), .C(n5461), .Y(n3459) );
  OAI21X1 U2720 ( .A(n10726), .B(n10781), .C(n5580), .Y(n3460) );
  OAI21X1 U2722 ( .A(n10726), .B(n10780), .C(n5696), .Y(n3461) );
  OAI21X1 U2724 ( .A(n10726), .B(n10779), .C(n4320), .Y(n3462) );
  OAI21X1 U2726 ( .A(n10725), .B(n10778), .C(n4319), .Y(n3463) );
  OAI21X1 U2728 ( .A(n10725), .B(n10777), .C(n5579), .Y(n3464) );
  OAI21X1 U2730 ( .A(n10725), .B(n10776), .C(n4318), .Y(n3465) );
  OAI21X1 U2732 ( .A(n10726), .B(n10775), .C(n4317), .Y(n3466) );
  OAI21X1 U2734 ( .A(n10726), .B(n10774), .C(n6088), .Y(n3467) );
  OAI21X1 U2736 ( .A(n10725), .B(n10773), .C(n5342), .Y(n3468) );
  OAI21X1 U2738 ( .A(n10726), .B(n10772), .C(n5460), .Y(n3469) );
  OAI21X1 U2740 ( .A(n10725), .B(n10771), .C(n6220), .Y(n3470) );
  OAI21X1 U2742 ( .A(n10725), .B(n10770), .C(n4316), .Y(n3471) );
  OAI21X1 U2744 ( .A(n10725), .B(n10769), .C(n5578), .Y(n3472) );
  OAI21X1 U2746 ( .A(n10726), .B(n10768), .C(n4315), .Y(n3473) );
  OAI21X1 U2748 ( .A(n10726), .B(n10767), .C(n5956), .Y(n3474) );
  OAI21X1 U2750 ( .A(n5653), .B(n6170), .C(reset_n), .Y(n1413) );
  OAI21X1 U2751 ( .A(n10723), .B(n10830), .C(n6219), .Y(n3475) );
  OAI21X1 U2753 ( .A(n10723), .B(n10829), .C(n6218), .Y(n3476) );
  OAI21X1 U2755 ( .A(n10723), .B(n10828), .C(n6087), .Y(n3477) );
  OAI21X1 U2757 ( .A(n10723), .B(n10827), .C(n5955), .Y(n3478) );
  OAI21X1 U2759 ( .A(n10723), .B(n10826), .C(n5823), .Y(n3479) );
  OAI21X1 U2761 ( .A(n10723), .B(n10825), .C(n5695), .Y(n3480) );
  OAI21X1 U2763 ( .A(n10723), .B(n10824), .C(n5577), .Y(n3481) );
  OAI21X1 U2765 ( .A(n10723), .B(n10823), .C(n5459), .Y(n3482) );
  OAI21X1 U2767 ( .A(n10723), .B(n10822), .C(n5341), .Y(n3483) );
  OAI21X1 U2769 ( .A(n10723), .B(n10821), .C(n5231), .Y(n3484) );
  OAI21X1 U2771 ( .A(n10723), .B(n10820), .C(n5122), .Y(n3485) );
  OAI21X1 U2773 ( .A(n10723), .B(n10819), .C(n5013), .Y(n3486) );
  OAI21X1 U2775 ( .A(n10723), .B(n10818), .C(n4904), .Y(n3487) );
  OAI21X1 U2777 ( .A(n10723), .B(n10817), .C(n6217), .Y(n3488) );
  OAI21X1 U2779 ( .A(n10723), .B(n10816), .C(n6086), .Y(n3489) );
  OAI21X1 U2781 ( .A(n10723), .B(n10815), .C(n5954), .Y(n3490) );
  OAI21X1 U2783 ( .A(n10724), .B(n10814), .C(n5822), .Y(n3491) );
  OAI21X1 U2785 ( .A(n10724), .B(n10813), .C(n5694), .Y(n3492) );
  OAI21X1 U2787 ( .A(n10723), .B(n10812), .C(n5576), .Y(n3493) );
  OAI21X1 U2789 ( .A(n10724), .B(n10811), .C(n5458), .Y(n3494) );
  OAI21X1 U2791 ( .A(n10724), .B(n10810), .C(n5340), .Y(n3495) );
  OAI21X1 U2793 ( .A(n10724), .B(n10809), .C(n5230), .Y(n3496) );
  OAI21X1 U2795 ( .A(n10724), .B(n10808), .C(n5121), .Y(n3497) );
  OAI21X1 U2797 ( .A(n10723), .B(n10807), .C(n5012), .Y(n3498) );
  OAI21X1 U2799 ( .A(n10723), .B(n10806), .C(n4796), .Y(n3499) );
  OAI21X1 U2801 ( .A(n10723), .B(n10805), .C(n5339), .Y(n3500) );
  OAI21X1 U2803 ( .A(n10723), .B(n10804), .C(n6085), .Y(n3501) );
  OAI21X1 U2805 ( .A(n10723), .B(n10803), .C(n5953), .Y(n3502) );
  OAI21X1 U2807 ( .A(n10724), .B(n10802), .C(n5821), .Y(n3503) );
  OAI21X1 U2809 ( .A(n10723), .B(n10801), .C(n5693), .Y(n3504) );
  OAI21X1 U2811 ( .A(n10724), .B(n10800), .C(n5575), .Y(n3505) );
  OAI21X1 U2813 ( .A(n10723), .B(n10799), .C(n5457), .Y(n3506) );
  OAI21X1 U2815 ( .A(n10723), .B(n10798), .C(n6216), .Y(n3507) );
  OAI21X1 U2817 ( .A(n10723), .B(n10797), .C(n5229), .Y(n3508) );
  OAI21X1 U2819 ( .A(n10724), .B(n10796), .C(n5120), .Y(n3509) );
  OAI21X1 U2821 ( .A(n10723), .B(n10795), .C(n5011), .Y(n3510) );
  OAI21X1 U2823 ( .A(n10723), .B(n10794), .C(n4903), .Y(n3511) );
  OAI21X1 U2825 ( .A(n10724), .B(n10793), .C(n6084), .Y(n3512) );
  OAI21X1 U2827 ( .A(n10723), .B(n10792), .C(n5574), .Y(n3513) );
  OAI21X1 U2829 ( .A(n10723), .B(n10791), .C(n5952), .Y(n3514) );
  OAI21X1 U2831 ( .A(n10723), .B(n10790), .C(n5820), .Y(n3515) );
  OAI21X1 U2833 ( .A(n10724), .B(n10789), .C(n5692), .Y(n3516) );
  OAI21X1 U2835 ( .A(n10724), .B(n10788), .C(n4902), .Y(n3517) );
  OAI21X1 U2837 ( .A(n10723), .B(n10787), .C(n5456), .Y(n3518) );
  OAI21X1 U2839 ( .A(n10724), .B(n10786), .C(n5228), .Y(n3519) );
  OAI21X1 U2841 ( .A(n10724), .B(n10785), .C(n6215), .Y(n3520) );
  OAI21X1 U2843 ( .A(n10723), .B(n10784), .C(n4795), .Y(n3521) );
  OAI21X1 U2845 ( .A(n10723), .B(n10783), .C(n5338), .Y(n3522) );
  OAI21X1 U2847 ( .A(n10723), .B(n10782), .C(n4689), .Y(n3523) );
  OAI21X1 U2849 ( .A(n10724), .B(n10781), .C(n4582), .Y(n3524) );
  OAI21X1 U2851 ( .A(n10724), .B(n10780), .C(n4475), .Y(n3525) );
  OAI21X1 U2853 ( .A(n10723), .B(n10779), .C(n4314), .Y(n3526) );
  OAI21X1 U2855 ( .A(n10724), .B(n10778), .C(n4313), .Y(n3527) );
  OAI21X1 U2857 ( .A(n10724), .B(n10777), .C(n4581), .Y(n3528) );
  OAI21X1 U2859 ( .A(n10723), .B(n10776), .C(n4312), .Y(n3529) );
  OAI21X1 U2861 ( .A(n10724), .B(n10775), .C(n4311), .Y(n3530) );
  OAI21X1 U2863 ( .A(n10724), .B(n10774), .C(n5010), .Y(n3531) );
  OAI21X1 U2865 ( .A(n10723), .B(n10773), .C(n4794), .Y(n3532) );
  OAI21X1 U2867 ( .A(n10724), .B(n10772), .C(n4688), .Y(n3533) );
  OAI21X1 U2869 ( .A(n10723), .B(n10771), .C(n4901), .Y(n3534) );
  OAI21X1 U2871 ( .A(n10723), .B(n10770), .C(n4310), .Y(n3535) );
  OAI21X1 U2873 ( .A(n10723), .B(n10769), .C(n4580), .Y(n3536) );
  OAI21X1 U2875 ( .A(n10724), .B(n10768), .C(n4309), .Y(n3537) );
  OAI21X1 U2877 ( .A(n10724), .B(n10767), .C(n5119), .Y(n3538) );
  OAI21X1 U2879 ( .A(n5771), .B(n6170), .C(reset_n), .Y(n1478) );
  OAI21X1 U2880 ( .A(n10721), .B(n10830), .C(n6083), .Y(n3539) );
  OAI21X1 U2882 ( .A(n10721), .B(n10829), .C(n6082), .Y(n3540) );
  OAI21X1 U2884 ( .A(n10721), .B(n10828), .C(n6214), .Y(n3541) );
  OAI21X1 U2886 ( .A(n10721), .B(n10827), .C(n5819), .Y(n3542) );
  OAI21X1 U2888 ( .A(n10721), .B(n10826), .C(n5951), .Y(n3543) );
  OAI21X1 U2890 ( .A(n10721), .B(n10825), .C(n5573), .Y(n3544) );
  OAI21X1 U2892 ( .A(n10721), .B(n10824), .C(n5691), .Y(n3545) );
  OAI21X1 U2894 ( .A(n10721), .B(n10823), .C(n5337), .Y(n3546) );
  OAI21X1 U2896 ( .A(n10721), .B(n10822), .C(n5455), .Y(n3547) );
  OAI21X1 U2898 ( .A(n10721), .B(n10821), .C(n5118), .Y(n3548) );
  OAI21X1 U2900 ( .A(n10721), .B(n10820), .C(n5227), .Y(n3549) );
  OAI21X1 U2902 ( .A(n10721), .B(n10819), .C(n4900), .Y(n3550) );
  OAI21X1 U2904 ( .A(n10721), .B(n10818), .C(n5009), .Y(n3551) );
  OAI21X1 U2906 ( .A(n10721), .B(n10817), .C(n6081), .Y(n3552) );
  OAI21X1 U2908 ( .A(n10721), .B(n10816), .C(n6213), .Y(n3553) );
  OAI21X1 U2910 ( .A(n10721), .B(n10815), .C(n5818), .Y(n3554) );
  OAI21X1 U2912 ( .A(n10722), .B(n10814), .C(n5950), .Y(n3555) );
  OAI21X1 U2914 ( .A(n10722), .B(n10813), .C(n5572), .Y(n3556) );
  OAI21X1 U2916 ( .A(n10721), .B(n10812), .C(n5690), .Y(n3557) );
  OAI21X1 U2918 ( .A(n10722), .B(n10811), .C(n5336), .Y(n3558) );
  OAI21X1 U2920 ( .A(n10722), .B(n10810), .C(n5454), .Y(n3559) );
  OAI21X1 U2922 ( .A(n10722), .B(n10809), .C(n5117), .Y(n3560) );
  OAI21X1 U2924 ( .A(n10722), .B(n10808), .C(n5226), .Y(n3561) );
  OAI21X1 U2926 ( .A(n10721), .B(n10807), .C(n4899), .Y(n3562) );
  OAI21X1 U2928 ( .A(n10721), .B(n10806), .C(n4687), .Y(n3563) );
  OAI21X1 U2930 ( .A(n10721), .B(n10805), .C(n5453), .Y(n3564) );
  OAI21X1 U2932 ( .A(n10721), .B(n10804), .C(n6212), .Y(n3565) );
  OAI21X1 U2934 ( .A(n10721), .B(n10803), .C(n5817), .Y(n3566) );
  OAI21X1 U2936 ( .A(n10722), .B(n10802), .C(n5949), .Y(n3567) );
  OAI21X1 U2938 ( .A(n10721), .B(n10801), .C(n5571), .Y(n3568) );
  OAI21X1 U2940 ( .A(n10722), .B(n10800), .C(n5689), .Y(n3569) );
  OAI21X1 U2942 ( .A(n10721), .B(n10799), .C(n5335), .Y(n3570) );
  OAI21X1 U2944 ( .A(n10721), .B(n10798), .C(n6080), .Y(n3571) );
  OAI21X1 U2946 ( .A(n10721), .B(n10797), .C(n5116), .Y(n3572) );
  OAI21X1 U2948 ( .A(n10722), .B(n10796), .C(n5225), .Y(n3573) );
  OAI21X1 U2950 ( .A(n10721), .B(n10795), .C(n4898), .Y(n3574) );
  OAI21X1 U2952 ( .A(n10721), .B(n10794), .C(n5008), .Y(n3575) );
  OAI21X1 U2954 ( .A(n10722), .B(n10793), .C(n6211), .Y(n3576) );
  OAI21X1 U2956 ( .A(n10721), .B(n10792), .C(n5688), .Y(n3577) );
  OAI21X1 U2958 ( .A(n10721), .B(n10791), .C(n5816), .Y(n3578) );
  OAI21X1 U2960 ( .A(n10721), .B(n10790), .C(n5948), .Y(n3579) );
  OAI21X1 U2962 ( .A(n10722), .B(n10789), .C(n5570), .Y(n3580) );
  OAI21X1 U2964 ( .A(n10722), .B(n10788), .C(n5007), .Y(n3581) );
  OAI21X1 U2966 ( .A(n10721), .B(n10787), .C(n5334), .Y(n3582) );
  OAI21X1 U2968 ( .A(n10722), .B(n10786), .C(n5115), .Y(n3583) );
  OAI21X1 U2970 ( .A(n10722), .B(n10785), .C(n6079), .Y(n3584) );
  OAI21X1 U2972 ( .A(n10721), .B(n10784), .C(n4686), .Y(n3585) );
  OAI21X1 U2974 ( .A(n10721), .B(n10783), .C(n5452), .Y(n3586) );
  OAI21X1 U2976 ( .A(n10721), .B(n10782), .C(n4793), .Y(n3587) );
  OAI21X1 U2978 ( .A(n10722), .B(n10781), .C(n4474), .Y(n3588) );
  OAI21X1 U2980 ( .A(n10722), .B(n10780), .C(n4579), .Y(n3589) );
  OAI21X1 U2982 ( .A(n10721), .B(n10779), .C(n4308), .Y(n3590) );
  OAI21X1 U2984 ( .A(n10722), .B(n10778), .C(n4307), .Y(n3591) );
  OAI21X1 U2986 ( .A(n10722), .B(n10777), .C(n4473), .Y(n3592) );
  OAI21X1 U2988 ( .A(n10721), .B(n10776), .C(n4306), .Y(n3593) );
  OAI21X1 U2990 ( .A(n10722), .B(n10775), .C(n4305), .Y(n3594) );
  OAI21X1 U2992 ( .A(n10722), .B(n10774), .C(n4897), .Y(n3595) );
  OAI21X1 U2994 ( .A(n10721), .B(n10773), .C(n4685), .Y(n3596) );
  OAI21X1 U2996 ( .A(n10722), .B(n10772), .C(n4792), .Y(n3597) );
  OAI21X1 U2998 ( .A(n10721), .B(n10771), .C(n5006), .Y(n3598) );
  OAI21X1 U3000 ( .A(n10721), .B(n10770), .C(n4304), .Y(n3599) );
  OAI21X1 U3002 ( .A(n10721), .B(n10769), .C(n4472), .Y(n3600) );
  OAI21X1 U3004 ( .A(n10722), .B(n10768), .C(n4303), .Y(n3601) );
  OAI21X1 U3006 ( .A(n10722), .B(n10767), .C(n5224), .Y(n3602) );
  OAI21X1 U3008 ( .A(n5535), .B(n6170), .C(reset_n), .Y(n1543) );
  OAI21X1 U3009 ( .A(n10719), .B(n10830), .C(n5947), .Y(n3603) );
  OAI21X1 U3011 ( .A(n10719), .B(n10829), .C(n5946), .Y(n3604) );
  OAI21X1 U3013 ( .A(n10719), .B(n10828), .C(n5815), .Y(n3605) );
  OAI21X1 U3015 ( .A(n10719), .B(n10827), .C(n6210), .Y(n3606) );
  OAI21X1 U3017 ( .A(n10719), .B(n10826), .C(n6078), .Y(n3607) );
  OAI21X1 U3019 ( .A(n10719), .B(n10825), .C(n5451), .Y(n3608) );
  OAI21X1 U3021 ( .A(n10719), .B(n10824), .C(n5333), .Y(n3609) );
  OAI21X1 U3023 ( .A(n10719), .B(n10823), .C(n5687), .Y(n3610) );
  OAI21X1 U3025 ( .A(n10719), .B(n10822), .C(n5569), .Y(n3611) );
  OAI21X1 U3027 ( .A(n10719), .B(n10821), .C(n5005), .Y(n3612) );
  OAI21X1 U3029 ( .A(n10719), .B(n10820), .C(n4896), .Y(n3613) );
  OAI21X1 U3031 ( .A(n10719), .B(n10819), .C(n5223), .Y(n3614) );
  OAI21X1 U3033 ( .A(n10719), .B(n10818), .C(n5114), .Y(n3615) );
  OAI21X1 U3035 ( .A(n10719), .B(n10817), .C(n5945), .Y(n3616) );
  OAI21X1 U3037 ( .A(n10719), .B(n10816), .C(n5814), .Y(n3617) );
  OAI21X1 U3039 ( .A(n10719), .B(n10815), .C(n6209), .Y(n3618) );
  OAI21X1 U3041 ( .A(n10720), .B(n10814), .C(n6077), .Y(n3619) );
  OAI21X1 U3043 ( .A(n10720), .B(n10813), .C(n5450), .Y(n3620) );
  OAI21X1 U3045 ( .A(n10719), .B(n10812), .C(n5332), .Y(n3621) );
  OAI21X1 U3047 ( .A(n10720), .B(n10811), .C(n5686), .Y(n3622) );
  OAI21X1 U3049 ( .A(n10720), .B(n10810), .C(n5568), .Y(n3623) );
  OAI21X1 U3051 ( .A(n10720), .B(n10809), .C(n5004), .Y(n3624) );
  OAI21X1 U3053 ( .A(n10720), .B(n10808), .C(n4895), .Y(n3625) );
  OAI21X1 U3055 ( .A(n10719), .B(n10807), .C(n5222), .Y(n3626) );
  OAI21X1 U3057 ( .A(n10719), .B(n10806), .C(n4578), .Y(n3627) );
  OAI21X1 U3059 ( .A(n10719), .B(n10805), .C(n5567), .Y(n3628) );
  OAI21X1 U3061 ( .A(n10719), .B(n10804), .C(n5813), .Y(n3629) );
  OAI21X1 U3063 ( .A(n10719), .B(n10803), .C(n6208), .Y(n3630) );
  OAI21X1 U3065 ( .A(n10720), .B(n10802), .C(n6076), .Y(n3631) );
  OAI21X1 U3067 ( .A(n10719), .B(n10801), .C(n5449), .Y(n3632) );
  OAI21X1 U3069 ( .A(n10720), .B(n10800), .C(n5331), .Y(n3633) );
  OAI21X1 U3071 ( .A(n10719), .B(n10799), .C(n5685), .Y(n3634) );
  OAI21X1 U3073 ( .A(n10719), .B(n10798), .C(n5944), .Y(n3635) );
  OAI21X1 U3075 ( .A(n10719), .B(n10797), .C(n5003), .Y(n3636) );
  OAI21X1 U3077 ( .A(n10720), .B(n10796), .C(n4894), .Y(n3637) );
  OAI21X1 U3079 ( .A(n10719), .B(n10795), .C(n5221), .Y(n3638) );
  OAI21X1 U3081 ( .A(n10719), .B(n10794), .C(n5113), .Y(n3639) );
  OAI21X1 U3083 ( .A(n10720), .B(n10793), .C(n5812), .Y(n3640) );
  OAI21X1 U3085 ( .A(n10719), .B(n10792), .C(n5330), .Y(n3641) );
  OAI21X1 U3087 ( .A(n10719), .B(n10791), .C(n6207), .Y(n3642) );
  OAI21X1 U3089 ( .A(n10719), .B(n10790), .C(n6075), .Y(n3643) );
  OAI21X1 U3091 ( .A(n10720), .B(n10789), .C(n5448), .Y(n3644) );
  OAI21X1 U3093 ( .A(n10720), .B(n10788), .C(n5112), .Y(n3645) );
  OAI21X1 U3095 ( .A(n10719), .B(n10787), .C(n5684), .Y(n3646) );
  OAI21X1 U3097 ( .A(n10720), .B(n10786), .C(n5002), .Y(n3647) );
  OAI21X1 U3099 ( .A(n10720), .B(n10785), .C(n5943), .Y(n3648) );
  OAI21X1 U3101 ( .A(n10719), .B(n10784), .C(n4577), .Y(n3649) );
  OAI21X1 U3103 ( .A(n10719), .B(n10783), .C(n5566), .Y(n3650) );
  OAI21X1 U3105 ( .A(n10719), .B(n10782), .C(n4471), .Y(n3651) );
  OAI21X1 U3107 ( .A(n10720), .B(n10781), .C(n4791), .Y(n3652) );
  OAI21X1 U3109 ( .A(n10720), .B(n10780), .C(n4684), .Y(n3653) );
  OAI21X1 U3111 ( .A(n10719), .B(n10779), .C(n4302), .Y(n3654) );
  OAI21X1 U3113 ( .A(n10720), .B(n10778), .C(n4301), .Y(n3655) );
  OAI21X1 U3115 ( .A(n10720), .B(n10777), .C(n4790), .Y(n3656) );
  OAI21X1 U3117 ( .A(n10719), .B(n10776), .C(n4300), .Y(n3657) );
  OAI21X1 U3119 ( .A(n10720), .B(n10775), .C(n4299), .Y(n3658) );
  OAI21X1 U3121 ( .A(n10720), .B(n10774), .C(n5220), .Y(n3659) );
  OAI21X1 U3123 ( .A(n10719), .B(n10773), .C(n4576), .Y(n3660) );
  OAI21X1 U3125 ( .A(n10720), .B(n10772), .C(n4470), .Y(n3661) );
  OAI21X1 U3127 ( .A(n10719), .B(n10771), .C(n5111), .Y(n3662) );
  OAI21X1 U3129 ( .A(n10719), .B(n10770), .C(n4298), .Y(n3663) );
  OAI21X1 U3131 ( .A(n10719), .B(n10769), .C(n4789), .Y(n3664) );
  OAI21X1 U3133 ( .A(n10720), .B(n10768), .C(n4297), .Y(n3665) );
  OAI21X1 U3135 ( .A(n10720), .B(n10767), .C(n4893), .Y(n3666) );
  OAI21X1 U3137 ( .A(n5417), .B(n6170), .C(reset_n), .Y(n1608) );
  OAI21X1 U3138 ( .A(n10717), .B(n10830), .C(n5811), .Y(n3667) );
  OAI21X1 U3140 ( .A(n10717), .B(n10829), .C(n5810), .Y(n3668) );
  OAI21X1 U3142 ( .A(n10717), .B(n10828), .C(n5942), .Y(n3669) );
  OAI21X1 U3144 ( .A(n10717), .B(n10827), .C(n6074), .Y(n3670) );
  OAI21X1 U3146 ( .A(n10717), .B(n10826), .C(n6206), .Y(n3671) );
  OAI21X1 U3148 ( .A(n10717), .B(n10825), .C(n5329), .Y(n3672) );
  OAI21X1 U3150 ( .A(n10717), .B(n10824), .C(n5447), .Y(n3673) );
  OAI21X1 U3152 ( .A(n10717), .B(n10823), .C(n5565), .Y(n3674) );
  OAI21X1 U3154 ( .A(n10717), .B(n10822), .C(n5683), .Y(n3675) );
  OAI21X1 U3156 ( .A(n10717), .B(n10821), .C(n4892), .Y(n3676) );
  OAI21X1 U3158 ( .A(n10717), .B(n10820), .C(n5001), .Y(n3677) );
  OAI21X1 U3160 ( .A(n10717), .B(n10819), .C(n5110), .Y(n3678) );
  OAI21X1 U3162 ( .A(n10717), .B(n10818), .C(n5219), .Y(n3679) );
  OAI21X1 U3164 ( .A(n10717), .B(n10817), .C(n5809), .Y(n3680) );
  OAI21X1 U3166 ( .A(n10717), .B(n10816), .C(n5941), .Y(n3681) );
  OAI21X1 U3168 ( .A(n10717), .B(n10815), .C(n6073), .Y(n3682) );
  OAI21X1 U3170 ( .A(n10718), .B(n10814), .C(n6205), .Y(n3683) );
  OAI21X1 U3172 ( .A(n10718), .B(n10813), .C(n5328), .Y(n3684) );
  OAI21X1 U3174 ( .A(n10717), .B(n10812), .C(n5446), .Y(n3685) );
  OAI21X1 U3176 ( .A(n10718), .B(n10811), .C(n5564), .Y(n3686) );
  OAI21X1 U3178 ( .A(n10718), .B(n10810), .C(n5682), .Y(n3687) );
  OAI21X1 U3180 ( .A(n10718), .B(n10809), .C(n4891), .Y(n3688) );
  OAI21X1 U3182 ( .A(n10718), .B(n10808), .C(n5000), .Y(n3689) );
  OAI21X1 U3184 ( .A(n10717), .B(n10807), .C(n5109), .Y(n3690) );
  OAI21X1 U3186 ( .A(n10717), .B(n10806), .C(n4469), .Y(n3691) );
  OAI21X1 U3188 ( .A(n10717), .B(n10805), .C(n5681), .Y(n3692) );
  OAI21X1 U3190 ( .A(n10717), .B(n10804), .C(n5940), .Y(n3693) );
  OAI21X1 U3192 ( .A(n10717), .B(n10803), .C(n6072), .Y(n3694) );
  OAI21X1 U3194 ( .A(n10718), .B(n10802), .C(n6204), .Y(n3695) );
  OAI21X1 U3196 ( .A(n10717), .B(n10801), .C(n5327), .Y(n3696) );
  OAI21X1 U3198 ( .A(n10718), .B(n10800), .C(n5445), .Y(n3697) );
  OAI21X1 U3200 ( .A(n10717), .B(n10799), .C(n5563), .Y(n3698) );
  OAI21X1 U3202 ( .A(n10717), .B(n10798), .C(n5808), .Y(n3699) );
  OAI21X1 U3204 ( .A(n10717), .B(n10797), .C(n4890), .Y(n3700) );
  OAI21X1 U3206 ( .A(n10718), .B(n10796), .C(n4999), .Y(n3701) );
  OAI21X1 U3208 ( .A(n10717), .B(n10795), .C(n5108), .Y(n3702) );
  OAI21X1 U3210 ( .A(n10717), .B(n10794), .C(n5218), .Y(n3703) );
  OAI21X1 U3212 ( .A(n10718), .B(n10793), .C(n5939), .Y(n3704) );
  OAI21X1 U3214 ( .A(n10717), .B(n10792), .C(n5444), .Y(n3705) );
  OAI21X1 U3216 ( .A(n10717), .B(n10791), .C(n6071), .Y(n3706) );
  OAI21X1 U3218 ( .A(n10717), .B(n10790), .C(n6203), .Y(n3707) );
  OAI21X1 U3220 ( .A(n10718), .B(n10789), .C(n5326), .Y(n3708) );
  OAI21X1 U3222 ( .A(n10718), .B(n10788), .C(n5217), .Y(n3709) );
  OAI21X1 U3224 ( .A(n10717), .B(n10787), .C(n5562), .Y(n3710) );
  OAI21X1 U3226 ( .A(n10718), .B(n10786), .C(n4889), .Y(n3711) );
  OAI21X1 U3228 ( .A(n10718), .B(n10785), .C(n5807), .Y(n3712) );
  OAI21X1 U3230 ( .A(n10717), .B(n10784), .C(n4468), .Y(n3713) );
  OAI21X1 U3232 ( .A(n10717), .B(n10783), .C(n5680), .Y(n3714) );
  OAI21X1 U3234 ( .A(n10717), .B(n10782), .C(n4575), .Y(n3715) );
  OAI21X1 U3236 ( .A(n10718), .B(n10781), .C(n4683), .Y(n3716) );
  OAI21X1 U3238 ( .A(n10718), .B(n10780), .C(n4788), .Y(n3717) );
  OAI21X1 U3240 ( .A(n10717), .B(n10779), .C(n4296), .Y(n3718) );
  OAI21X1 U3242 ( .A(n10718), .B(n10778), .C(n4295), .Y(n3719) );
  OAI21X1 U3244 ( .A(n10718), .B(n10777), .C(n4682), .Y(n3720) );
  OAI21X1 U3246 ( .A(n10717), .B(n10776), .C(n4294), .Y(n3721) );
  OAI21X1 U3248 ( .A(n10718), .B(n10775), .C(n4293), .Y(n3722) );
  OAI21X1 U3250 ( .A(n10718), .B(n10774), .C(n5107), .Y(n3723) );
  OAI21X1 U3252 ( .A(n10717), .B(n10773), .C(n4467), .Y(n3724) );
  OAI21X1 U3254 ( .A(n10718), .B(n10772), .C(n4574), .Y(n3725) );
  OAI21X1 U3256 ( .A(n10717), .B(n10771), .C(n5216), .Y(n3726) );
  OAI21X1 U3258 ( .A(n10717), .B(n10770), .C(n4292), .Y(n3727) );
  OAI21X1 U3260 ( .A(n10717), .B(n10769), .C(n4681), .Y(n3728) );
  OAI21X1 U3262 ( .A(n10718), .B(n10768), .C(n4291), .Y(n3729) );
  OAI21X1 U3264 ( .A(n10718), .B(n10767), .C(n4998), .Y(n3730) );
  OAI21X1 U3266 ( .A(n5299), .B(n6170), .C(reset_n), .Y(n1673) );
  NAND3X1 U3267 ( .A(n10765), .B(n10831), .C(waddr[3]), .Y(n1218) );
  OAI21X1 U3268 ( .A(n10715), .B(n10830), .C(n5679), .Y(n3731) );
  OAI21X1 U3270 ( .A(n10715), .B(n10829), .C(n5678), .Y(n3732) );
  OAI21X1 U3272 ( .A(n10715), .B(n10828), .C(n5561), .Y(n3733) );
  OAI21X1 U3274 ( .A(n10715), .B(n10827), .C(n5443), .Y(n3734) );
  OAI21X1 U3276 ( .A(n10715), .B(n10826), .C(n5325), .Y(n3735) );
  OAI21X1 U3278 ( .A(n10715), .B(n10825), .C(n6202), .Y(n3736) );
  OAI21X1 U3280 ( .A(n10715), .B(n10824), .C(n6070), .Y(n3737) );
  OAI21X1 U3282 ( .A(n10715), .B(n10823), .C(n5938), .Y(n3738) );
  OAI21X1 U3284 ( .A(n10715), .B(n10822), .C(n5806), .Y(n3739) );
  OAI21X1 U3286 ( .A(n10715), .B(n10821), .C(n4787), .Y(n3740) );
  OAI21X1 U3288 ( .A(n10715), .B(n10820), .C(n4680), .Y(n3741) );
  OAI21X1 U3290 ( .A(n10715), .B(n10819), .C(n4573), .Y(n3742) );
  OAI21X1 U3292 ( .A(n10715), .B(n10818), .C(n4466), .Y(n3743) );
  OAI21X1 U3294 ( .A(n10715), .B(n10817), .C(n5677), .Y(n3744) );
  OAI21X1 U3296 ( .A(n10715), .B(n10816), .C(n5560), .Y(n3745) );
  OAI21X1 U3298 ( .A(n10715), .B(n10815), .C(n5442), .Y(n3746) );
  OAI21X1 U3300 ( .A(n10716), .B(n10814), .C(n5324), .Y(n3747) );
  OAI21X1 U3302 ( .A(n10716), .B(n10813), .C(n6201), .Y(n3748) );
  OAI21X1 U3304 ( .A(n10715), .B(n10812), .C(n6069), .Y(n3749) );
  OAI21X1 U3306 ( .A(n10716), .B(n10811), .C(n5937), .Y(n3750) );
  OAI21X1 U3308 ( .A(n10716), .B(n10810), .C(n5805), .Y(n3751) );
  OAI21X1 U3310 ( .A(n10716), .B(n10809), .C(n4786), .Y(n3752) );
  OAI21X1 U3312 ( .A(n10716), .B(n10808), .C(n4679), .Y(n3753) );
  OAI21X1 U3314 ( .A(n10715), .B(n10807), .C(n4572), .Y(n3754) );
  OAI21X1 U3316 ( .A(n10715), .B(n10806), .C(n5215), .Y(n3755) );
  OAI21X1 U3318 ( .A(n10715), .B(n10805), .C(n5804), .Y(n3756) );
  OAI21X1 U3320 ( .A(n10715), .B(n10804), .C(n5559), .Y(n3757) );
  OAI21X1 U3322 ( .A(n10715), .B(n10803), .C(n5441), .Y(n3758) );
  OAI21X1 U3324 ( .A(n10716), .B(n10802), .C(n5323), .Y(n3759) );
  OAI21X1 U3326 ( .A(n10715), .B(n10801), .C(n6200), .Y(n3760) );
  OAI21X1 U3328 ( .A(n10716), .B(n10800), .C(n6068), .Y(n3761) );
  OAI21X1 U3330 ( .A(n10715), .B(n10799), .C(n5936), .Y(n3762) );
  OAI21X1 U3332 ( .A(n10715), .B(n10798), .C(n5676), .Y(n3763) );
  OAI21X1 U3334 ( .A(n10715), .B(n10797), .C(n4785), .Y(n3764) );
  OAI21X1 U3336 ( .A(n10716), .B(n10796), .C(n4678), .Y(n3765) );
  OAI21X1 U3338 ( .A(n10715), .B(n10795), .C(n4571), .Y(n3766) );
  OAI21X1 U3340 ( .A(n10715), .B(n10794), .C(n4465), .Y(n3767) );
  OAI21X1 U3342 ( .A(n10716), .B(n10793), .C(n5558), .Y(n3768) );
  OAI21X1 U3344 ( .A(n10715), .B(n10792), .C(n6067), .Y(n3769) );
  OAI21X1 U3346 ( .A(n10715), .B(n10791), .C(n5440), .Y(n3770) );
  OAI21X1 U3348 ( .A(n10715), .B(n10790), .C(n5322), .Y(n3771) );
  OAI21X1 U3350 ( .A(n10716), .B(n10789), .C(n6199), .Y(n3772) );
  OAI21X1 U3352 ( .A(n10716), .B(n10788), .C(n4464), .Y(n3773) );
  OAI21X1 U3354 ( .A(n10715), .B(n10787), .C(n5935), .Y(n3774) );
  OAI21X1 U3356 ( .A(n10716), .B(n10786), .C(n4784), .Y(n3775) );
  OAI21X1 U3358 ( .A(n10716), .B(n10785), .C(n5675), .Y(n3776) );
  OAI21X1 U3360 ( .A(n10715), .B(n10784), .C(n5214), .Y(n3777) );
  OAI21X1 U3362 ( .A(n10715), .B(n10783), .C(n5803), .Y(n3778) );
  OAI21X1 U3364 ( .A(n10715), .B(n10782), .C(n5106), .Y(n3779) );
  OAI21X1 U3366 ( .A(n10716), .B(n10781), .C(n4997), .Y(n3780) );
  OAI21X1 U3368 ( .A(n10716), .B(n10780), .C(n4888), .Y(n3781) );
  OAI21X1 U3370 ( .A(n10715), .B(n10779), .C(n4290), .Y(n3782) );
  OAI21X1 U3372 ( .A(n10716), .B(n10778), .C(n4289), .Y(n3783) );
  OAI21X1 U3374 ( .A(n10716), .B(n10777), .C(n4996), .Y(n3784) );
  OAI21X1 U3376 ( .A(n10715), .B(n10776), .C(n4288), .Y(n3785) );
  OAI21X1 U3378 ( .A(n10716), .B(n10775), .C(n4287), .Y(n3786) );
  OAI21X1 U3380 ( .A(n10716), .B(n10774), .C(n4570), .Y(n3787) );
  OAI21X1 U3382 ( .A(n10715), .B(n10773), .C(n5213), .Y(n3788) );
  OAI21X1 U3384 ( .A(n10716), .B(n10772), .C(n5105), .Y(n3789) );
  OAI21X1 U3386 ( .A(n10715), .B(n10771), .C(n4463), .Y(n3790) );
  OAI21X1 U3388 ( .A(n10715), .B(n10770), .C(n4286), .Y(n3791) );
  OAI21X1 U3390 ( .A(n10715), .B(n10769), .C(n4995), .Y(n3792) );
  OAI21X1 U3392 ( .A(n10716), .B(n10768), .C(n4285), .Y(n3793) );
  OAI21X1 U3394 ( .A(n10716), .B(n10767), .C(n4677), .Y(n3794) );
  OAI21X1 U3396 ( .A(n5774), .B(n6038), .C(reset_n), .Y(n1738) );
  NAND3X1 U3397 ( .A(waddr[1]), .B(waddr[0]), .C(waddr[2]), .Y(n168) );
  OAI21X1 U3398 ( .A(n10713), .B(n10830), .C(n5557), .Y(n3795) );
  OAI21X1 U3400 ( .A(n10713), .B(n10829), .C(n5556), .Y(n3796) );
  OAI21X1 U3402 ( .A(n10713), .B(n10828), .C(n5674), .Y(n3797) );
  OAI21X1 U3404 ( .A(n10713), .B(n10827), .C(n5321), .Y(n3798) );
  OAI21X1 U3406 ( .A(n10713), .B(n10826), .C(n5439), .Y(n3799) );
  OAI21X1 U3408 ( .A(n10713), .B(n10825), .C(n6066), .Y(n3800) );
  OAI21X1 U3410 ( .A(n10713), .B(n10824), .C(n6198), .Y(n3801) );
  OAI21X1 U3412 ( .A(n10713), .B(n10823), .C(n5802), .Y(n3802) );
  OAI21X1 U3414 ( .A(n10713), .B(n10822), .C(n5934), .Y(n3803) );
  OAI21X1 U3416 ( .A(n10713), .B(n10821), .C(n4676), .Y(n3804) );
  OAI21X1 U3418 ( .A(n10713), .B(n10820), .C(n4783), .Y(n3805) );
  OAI21X1 U3420 ( .A(n10713), .B(n10819), .C(n4462), .Y(n3806) );
  OAI21X1 U3422 ( .A(n10713), .B(n10818), .C(n4569), .Y(n3807) );
  OAI21X1 U3424 ( .A(n10713), .B(n10817), .C(n5555), .Y(n3808) );
  OAI21X1 U3426 ( .A(n10713), .B(n10816), .C(n5673), .Y(n3809) );
  OAI21X1 U3428 ( .A(n10713), .B(n10815), .C(n5320), .Y(n3810) );
  OAI21X1 U3430 ( .A(n10714), .B(n10814), .C(n5438), .Y(n3811) );
  OAI21X1 U3432 ( .A(n10714), .B(n10813), .C(n6065), .Y(n3812) );
  OAI21X1 U3434 ( .A(n10713), .B(n10812), .C(n6197), .Y(n3813) );
  OAI21X1 U3436 ( .A(n10714), .B(n10811), .C(n5801), .Y(n3814) );
  OAI21X1 U3438 ( .A(n10714), .B(n10810), .C(n5933), .Y(n3815) );
  OAI21X1 U3440 ( .A(n10714), .B(n10809), .C(n4675), .Y(n3816) );
  OAI21X1 U3442 ( .A(n10714), .B(n10808), .C(n4782), .Y(n3817) );
  OAI21X1 U3444 ( .A(n10713), .B(n10807), .C(n4461), .Y(n3818) );
  OAI21X1 U3446 ( .A(n10713), .B(n10806), .C(n5104), .Y(n3819) );
  OAI21X1 U3448 ( .A(n10713), .B(n10805), .C(n5932), .Y(n3820) );
  OAI21X1 U3450 ( .A(n10713), .B(n10804), .C(n5672), .Y(n3821) );
  OAI21X1 U3452 ( .A(n10713), .B(n10803), .C(n5319), .Y(n3822) );
  OAI21X1 U3454 ( .A(n10714), .B(n10802), .C(n5437), .Y(n3823) );
  OAI21X1 U3456 ( .A(n10713), .B(n10801), .C(n6064), .Y(n3824) );
  OAI21X1 U3458 ( .A(n10714), .B(n10800), .C(n6196), .Y(n3825) );
  OAI21X1 U3460 ( .A(n10713), .B(n10799), .C(n5800), .Y(n3826) );
  OAI21X1 U3462 ( .A(n10713), .B(n10798), .C(n5554), .Y(n3827) );
  OAI21X1 U3464 ( .A(n10713), .B(n10797), .C(n4674), .Y(n3828) );
  OAI21X1 U3466 ( .A(n10714), .B(n10796), .C(n4781), .Y(n3829) );
  OAI21X1 U3468 ( .A(n10713), .B(n10795), .C(n4460), .Y(n3830) );
  OAI21X1 U3470 ( .A(n10713), .B(n10794), .C(n4568), .Y(n3831) );
  OAI21X1 U3472 ( .A(n10714), .B(n10793), .C(n5671), .Y(n3832) );
  OAI21X1 U3474 ( .A(n10713), .B(n10792), .C(n6195), .Y(n3833) );
  OAI21X1 U3476 ( .A(n10713), .B(n10791), .C(n5318), .Y(n3834) );
  OAI21X1 U3478 ( .A(n10713), .B(n10790), .C(n5436), .Y(n3835) );
  OAI21X1 U3480 ( .A(n10714), .B(n10789), .C(n6063), .Y(n3836) );
  OAI21X1 U3482 ( .A(n10714), .B(n10788), .C(n4567), .Y(n3837) );
  OAI21X1 U3484 ( .A(n10713), .B(n10787), .C(n5799), .Y(n3838) );
  OAI21X1 U3486 ( .A(n10714), .B(n10786), .C(n4673), .Y(n3839) );
  OAI21X1 U3488 ( .A(n10714), .B(n10785), .C(n5553), .Y(n3840) );
  OAI21X1 U3490 ( .A(n10713), .B(n10784), .C(n5103), .Y(n3841) );
  OAI21X1 U3492 ( .A(n10713), .B(n10783), .C(n5931), .Y(n3842) );
  OAI21X1 U3494 ( .A(n10713), .B(n10782), .C(n5212), .Y(n3843) );
  OAI21X1 U3496 ( .A(n10714), .B(n10781), .C(n4887), .Y(n3844) );
  OAI21X1 U3498 ( .A(n10714), .B(n10780), .C(n4994), .Y(n3845) );
  OAI21X1 U3500 ( .A(n10713), .B(n10779), .C(n4284), .Y(n3846) );
  OAI21X1 U3502 ( .A(n10714), .B(n10778), .C(n4283), .Y(n3847) );
  OAI21X1 U3504 ( .A(n10714), .B(n10777), .C(n4886), .Y(n3848) );
  OAI21X1 U3506 ( .A(n10713), .B(n10776), .C(n4282), .Y(n3849) );
  OAI21X1 U3508 ( .A(n10714), .B(n10775), .C(n4281), .Y(n3850) );
  OAI21X1 U3510 ( .A(n10714), .B(n10774), .C(n4459), .Y(n3851) );
  OAI21X1 U3512 ( .A(n10713), .B(n10773), .C(n5102), .Y(n3852) );
  OAI21X1 U3514 ( .A(n10714), .B(n10772), .C(n5211), .Y(n3853) );
  OAI21X1 U3516 ( .A(n10713), .B(n10771), .C(n4566), .Y(n3854) );
  OAI21X1 U3518 ( .A(n10713), .B(n10770), .C(n4280), .Y(n3855) );
  OAI21X1 U3520 ( .A(n10713), .B(n10769), .C(n4885), .Y(n3856) );
  OAI21X1 U3522 ( .A(n10714), .B(n10768), .C(n4279), .Y(n3857) );
  OAI21X1 U3524 ( .A(n10714), .B(n10767), .C(n4780), .Y(n3858) );
  OAI21X1 U3526 ( .A(n5773), .B(n6038), .C(reset_n), .Y(n1804) );
  NAND3X1 U3527 ( .A(waddr[1]), .B(n10835), .C(waddr[2]), .Y(n234) );
  OAI21X1 U3528 ( .A(n10711), .B(n10830), .C(n5435), .Y(n3859) );
  OAI21X1 U3530 ( .A(n10711), .B(n10829), .C(n5434), .Y(n3860) );
  OAI21X1 U3532 ( .A(n10711), .B(n10828), .C(n5317), .Y(n3861) );
  OAI21X1 U3534 ( .A(n10711), .B(n10827), .C(n5670), .Y(n3862) );
  OAI21X1 U3536 ( .A(n10711), .B(n10826), .C(n5552), .Y(n3863) );
  OAI21X1 U3538 ( .A(n10711), .B(n10825), .C(n5930), .Y(n3864) );
  OAI21X1 U3540 ( .A(n10711), .B(n10824), .C(n5798), .Y(n3865) );
  OAI21X1 U3542 ( .A(n10711), .B(n10823), .C(n6194), .Y(n3866) );
  OAI21X1 U3544 ( .A(n10711), .B(n10822), .C(n6062), .Y(n3867) );
  OAI21X1 U3546 ( .A(n10711), .B(n10821), .C(n4565), .Y(n3868) );
  OAI21X1 U3548 ( .A(n10711), .B(n10820), .C(n4458), .Y(n3869) );
  OAI21X1 U3550 ( .A(n10711), .B(n10819), .C(n4779), .Y(n3870) );
  OAI21X1 U3552 ( .A(n10711), .B(n10818), .C(n4672), .Y(n3871) );
  OAI21X1 U3554 ( .A(n10711), .B(n10817), .C(n5433), .Y(n3872) );
  OAI21X1 U3556 ( .A(n10711), .B(n10816), .C(n5316), .Y(n3873) );
  OAI21X1 U3558 ( .A(n10711), .B(n10815), .C(n5669), .Y(n3874) );
  OAI21X1 U3560 ( .A(n10712), .B(n10814), .C(n5551), .Y(n3875) );
  OAI21X1 U3562 ( .A(n10712), .B(n10813), .C(n5929), .Y(n3876) );
  OAI21X1 U3564 ( .A(n10711), .B(n10812), .C(n5797), .Y(n3877) );
  OAI21X1 U3566 ( .A(n10712), .B(n10811), .C(n6193), .Y(n3878) );
  OAI21X1 U3568 ( .A(n10712), .B(n10810), .C(n6061), .Y(n3879) );
  OAI21X1 U3570 ( .A(n10712), .B(n10809), .C(n4564), .Y(n3880) );
  OAI21X1 U3572 ( .A(n10712), .B(n10808), .C(n4457), .Y(n3881) );
  OAI21X1 U3574 ( .A(n10711), .B(n10807), .C(n4778), .Y(n3882) );
  OAI21X1 U3576 ( .A(n10711), .B(n10806), .C(n4993), .Y(n3883) );
  OAI21X1 U3578 ( .A(n10711), .B(n10805), .C(n6060), .Y(n3884) );
  OAI21X1 U3580 ( .A(n10711), .B(n10804), .C(n5315), .Y(n3885) );
  OAI21X1 U3582 ( .A(n10711), .B(n10803), .C(n5668), .Y(n3886) );
  OAI21X1 U3584 ( .A(n10712), .B(n10802), .C(n5550), .Y(n3887) );
  OAI21X1 U3586 ( .A(n10711), .B(n10801), .C(n5928), .Y(n3888) );
  OAI21X1 U3588 ( .A(n10712), .B(n10800), .C(n5796), .Y(n3889) );
  OAI21X1 U3590 ( .A(n10711), .B(n10799), .C(n6192), .Y(n3890) );
  OAI21X1 U3592 ( .A(n10711), .B(n10798), .C(n5432), .Y(n3891) );
  OAI21X1 U3594 ( .A(n10711), .B(n10797), .C(n4563), .Y(n3892) );
  OAI21X1 U3596 ( .A(n10712), .B(n10796), .C(n4456), .Y(n3893) );
  OAI21X1 U3598 ( .A(n10711), .B(n10795), .C(n4777), .Y(n3894) );
  OAI21X1 U3600 ( .A(n10711), .B(n10794), .C(n4671), .Y(n3895) );
  OAI21X1 U3602 ( .A(n10712), .B(n10793), .C(n5314), .Y(n3896) );
  OAI21X1 U3604 ( .A(n10711), .B(n10792), .C(n5795), .Y(n3897) );
  OAI21X1 U3606 ( .A(n10711), .B(n10791), .C(n5667), .Y(n3898) );
  OAI21X1 U3608 ( .A(n10711), .B(n10790), .C(n5549), .Y(n3899) );
  OAI21X1 U3610 ( .A(n10712), .B(n10789), .C(n5927), .Y(n3900) );
  OAI21X1 U3612 ( .A(n10712), .B(n10788), .C(n4670), .Y(n3901) );
  OAI21X1 U3614 ( .A(n10711), .B(n10787), .C(n6191), .Y(n3902) );
  OAI21X1 U3616 ( .A(n10712), .B(n10786), .C(n4562), .Y(n3903) );
  OAI21X1 U3618 ( .A(n10712), .B(n10785), .C(n5431), .Y(n3904) );
  OAI21X1 U3620 ( .A(n10711), .B(n10784), .C(n4992), .Y(n3905) );
  OAI21X1 U3622 ( .A(n10711), .B(n10783), .C(n6059), .Y(n3906) );
  OAI21X1 U3624 ( .A(n10711), .B(n10782), .C(n4884), .Y(n3907) );
  OAI21X1 U3626 ( .A(n10712), .B(n10781), .C(n5210), .Y(n3908) );
  OAI21X1 U3628 ( .A(n10712), .B(n10780), .C(n5101), .Y(n3909) );
  OAI21X1 U3630 ( .A(n10711), .B(n10779), .C(n4278), .Y(n3910) );
  OAI21X1 U3632 ( .A(n10712), .B(n10778), .C(n4277), .Y(n3911) );
  OAI21X1 U3634 ( .A(n10712), .B(n10777), .C(n5209), .Y(n3912) );
  OAI21X1 U3636 ( .A(n10711), .B(n10776), .C(n4276), .Y(n3913) );
  OAI21X1 U3638 ( .A(n10712), .B(n10775), .C(n4275), .Y(n3914) );
  OAI21X1 U3640 ( .A(n10712), .B(n10774), .C(n4776), .Y(n3915) );
  OAI21X1 U3642 ( .A(n10711), .B(n10773), .C(n4991), .Y(n3916) );
  OAI21X1 U3644 ( .A(n10712), .B(n10772), .C(n4883), .Y(n3917) );
  OAI21X1 U3646 ( .A(n10711), .B(n10771), .C(n4669), .Y(n3918) );
  OAI21X1 U3648 ( .A(n10711), .B(n10770), .C(n4274), .Y(n3919) );
  OAI21X1 U3650 ( .A(n10711), .B(n10769), .C(n5208), .Y(n3920) );
  OAI21X1 U3652 ( .A(n10712), .B(n10768), .C(n4273), .Y(n3921) );
  OAI21X1 U3654 ( .A(n10712), .B(n10767), .C(n4455), .Y(n3922) );
  OAI21X1 U3656 ( .A(n5772), .B(n6038), .C(reset_n), .Y(n1869) );
  NAND3X1 U3657 ( .A(waddr[0]), .B(n10834), .C(waddr[2]), .Y(n300) );
  OAI21X1 U3658 ( .A(n10709), .B(n10830), .C(n5313), .Y(n3923) );
  OAI21X1 U3660 ( .A(n10709), .B(n10829), .C(n5312), .Y(n3924) );
  OAI21X1 U3662 ( .A(n10709), .B(n10828), .C(n5430), .Y(n3925) );
  OAI21X1 U3664 ( .A(n10709), .B(n10827), .C(n5548), .Y(n3926) );
  OAI21X1 U3666 ( .A(n10709), .B(n10826), .C(n5666), .Y(n3927) );
  OAI21X1 U3668 ( .A(n10709), .B(n10825), .C(n5794), .Y(n3928) );
  OAI21X1 U3670 ( .A(n10709), .B(n10824), .C(n5926), .Y(n3929) );
  OAI21X1 U3672 ( .A(n10709), .B(n10823), .C(n6058), .Y(n3930) );
  OAI21X1 U3674 ( .A(n10709), .B(n10822), .C(n6190), .Y(n3931) );
  OAI21X1 U3676 ( .A(n10709), .B(n10821), .C(n4454), .Y(n3932) );
  OAI21X1 U3678 ( .A(n10709), .B(n10820), .C(n4561), .Y(n3933) );
  OAI21X1 U3680 ( .A(n10709), .B(n10819), .C(n4668), .Y(n3934) );
  OAI21X1 U3682 ( .A(n10709), .B(n10818), .C(n4775), .Y(n3935) );
  OAI21X1 U3684 ( .A(n10709), .B(n10817), .C(n5311), .Y(n3936) );
  OAI21X1 U3686 ( .A(n10709), .B(n10816), .C(n5429), .Y(n3937) );
  OAI21X1 U3688 ( .A(n10710), .B(n10815), .C(n5547), .Y(n3938) );
  OAI21X1 U3690 ( .A(n10709), .B(n10814), .C(n5665), .Y(n3939) );
  OAI21X1 U3692 ( .A(n10710), .B(n10813), .C(n5793), .Y(n3940) );
  OAI21X1 U3694 ( .A(n10709), .B(n10812), .C(n5925), .Y(n3941) );
  OAI21X1 U3696 ( .A(n10710), .B(n10811), .C(n6057), .Y(n3942) );
  OAI21X1 U3698 ( .A(n10710), .B(n10810), .C(n6189), .Y(n3943) );
  OAI21X1 U3700 ( .A(n10710), .B(n10809), .C(n4453), .Y(n3944) );
  OAI21X1 U3702 ( .A(n10710), .B(n10808), .C(n4560), .Y(n3945) );
  OAI21X1 U3704 ( .A(n10709), .B(n10807), .C(n4667), .Y(n3946) );
  OAI21X1 U3706 ( .A(n10709), .B(n10806), .C(n4882), .Y(n3947) );
  OAI21X1 U3708 ( .A(n10709), .B(n10805), .C(n6188), .Y(n3948) );
  OAI21X1 U3710 ( .A(n10709), .B(n10804), .C(n5428), .Y(n3949) );
  OAI21X1 U3712 ( .A(n10709), .B(n10803), .C(n5546), .Y(n3950) );
  OAI21X1 U3714 ( .A(n10710), .B(n10802), .C(n5664), .Y(n3951) );
  OAI21X1 U3716 ( .A(n10710), .B(n10801), .C(n5792), .Y(n3952) );
  OAI21X1 U3718 ( .A(n10710), .B(n10800), .C(n5924), .Y(n3953) );
  OAI21X1 U3720 ( .A(n10709), .B(n10799), .C(n6056), .Y(n3954) );
  OAI21X1 U3722 ( .A(n10709), .B(n10798), .C(n5310), .Y(n3955) );
  OAI21X1 U3724 ( .A(n10709), .B(n10797), .C(n4452), .Y(n3956) );
  OAI21X1 U3726 ( .A(n10709), .B(n10796), .C(n4559), .Y(n3957) );
  OAI21X1 U3728 ( .A(n10710), .B(n10795), .C(n4666), .Y(n3958) );
  OAI21X1 U3730 ( .A(n10709), .B(n10794), .C(n4774), .Y(n3959) );
  OAI21X1 U3732 ( .A(n10709), .B(n10793), .C(n5427), .Y(n3960) );
  OAI21X1 U3734 ( .A(n10709), .B(n10792), .C(n5923), .Y(n3961) );
  OAI21X1 U3736 ( .A(n10709), .B(n10791), .C(n5545), .Y(n3962) );
  OAI21X1 U3738 ( .A(n10709), .B(n10790), .C(n5663), .Y(n3963) );
  OAI21X1 U3740 ( .A(n10710), .B(n10789), .C(n5791), .Y(n3964) );
  OAI21X1 U3742 ( .A(n10710), .B(n10788), .C(n4773), .Y(n3965) );
  OAI21X1 U3744 ( .A(n10709), .B(n10787), .C(n6055), .Y(n3966) );
  OAI21X1 U3746 ( .A(n10710), .B(n10786), .C(n4451), .Y(n3967) );
  OAI21X1 U3748 ( .A(n10710), .B(n10785), .C(n5309), .Y(n3968) );
  OAI21X1 U3750 ( .A(n10709), .B(n10784), .C(n4881), .Y(n3969) );
  OAI21X1 U3752 ( .A(n10710), .B(n10783), .C(n6187), .Y(n3970) );
  OAI21X1 U3754 ( .A(n10709), .B(n10782), .C(n4990), .Y(n3971) );
  OAI21X1 U3756 ( .A(n10710), .B(n10781), .C(n5100), .Y(n3972) );
  OAI21X1 U3758 ( .A(n10710), .B(n10780), .C(n5207), .Y(n3973) );
  OAI21X1 U3760 ( .A(n10710), .B(n10779), .C(n4272), .Y(n3974) );
  OAI21X1 U3762 ( .A(n10709), .B(n10778), .C(n4271), .Y(n3975) );
  OAI21X1 U3764 ( .A(n10709), .B(n10777), .C(n5099), .Y(n3976) );
  OAI21X1 U3766 ( .A(n10709), .B(n10776), .C(n4270), .Y(n3977) );
  OAI21X1 U3768 ( .A(n10710), .B(n10775), .C(n4269), .Y(n3978) );
  OAI21X1 U3770 ( .A(n10710), .B(n10774), .C(n4665), .Y(n3979) );
  OAI21X1 U3772 ( .A(n10709), .B(n10773), .C(n4880), .Y(n3980) );
  OAI21X1 U3774 ( .A(n10710), .B(n10772), .C(n4989), .Y(n3981) );
  OAI21X1 U3776 ( .A(n10709), .B(n10771), .C(n4772), .Y(n3982) );
  OAI21X1 U3778 ( .A(n10709), .B(n10770), .C(n4268), .Y(n3983) );
  OAI21X1 U3780 ( .A(n10709), .B(n10769), .C(n5098), .Y(n3984) );
  OAI21X1 U3782 ( .A(n10710), .B(n10768), .C(n4267), .Y(n3985) );
  OAI21X1 U3784 ( .A(n10710), .B(n10767), .C(n4558), .Y(n3986) );
  OAI21X1 U3786 ( .A(n5653), .B(n6038), .C(reset_n), .Y(n1934) );
  NAND3X1 U3787 ( .A(n10835), .B(n10834), .C(waddr[2]), .Y(n366) );
  OAI21X1 U3788 ( .A(n10707), .B(n10830), .C(n5206), .Y(n3987) );
  OAI21X1 U3790 ( .A(n10707), .B(n10829), .C(n5205), .Y(n3988) );
  OAI21X1 U3792 ( .A(n10707), .B(n10828), .C(n5097), .Y(n3989) );
  OAI21X1 U3794 ( .A(n10707), .B(n10827), .C(n4988), .Y(n3990) );
  OAI21X1 U3796 ( .A(n10707), .B(n10826), .C(n4879), .Y(n3991) );
  OAI21X1 U3798 ( .A(n10707), .B(n10825), .C(n4771), .Y(n3992) );
  OAI21X1 U3800 ( .A(n10707), .B(n10824), .C(n4664), .Y(n3993) );
  OAI21X1 U3802 ( .A(n10707), .B(n10823), .C(n4557), .Y(n3994) );
  OAI21X1 U3804 ( .A(n10707), .B(n10822), .C(n4450), .Y(n3995) );
  OAI21X1 U3806 ( .A(n10707), .B(n10821), .C(n6186), .Y(n3996) );
  OAI21X1 U3808 ( .A(n10707), .B(n10820), .C(n6054), .Y(n3997) );
  OAI21X1 U3810 ( .A(n10707), .B(n10819), .C(n5922), .Y(n3998) );
  OAI21X1 U3812 ( .A(n10707), .B(n10818), .C(n5790), .Y(n3999) );
  OAI21X1 U3814 ( .A(n10707), .B(n10817), .C(n5204), .Y(n4000) );
  OAI21X1 U3816 ( .A(n10707), .B(n10816), .C(n5096), .Y(n4001) );
  OAI21X1 U3818 ( .A(n10708), .B(n10815), .C(n4987), .Y(n4002) );
  OAI21X1 U3820 ( .A(n10707), .B(n10814), .C(n4878), .Y(n4003) );
  OAI21X1 U3822 ( .A(n10708), .B(n10813), .C(n4770), .Y(n4004) );
  OAI21X1 U3824 ( .A(n10707), .B(n10812), .C(n4663), .Y(n4005) );
  OAI21X1 U3826 ( .A(n10708), .B(n10811), .C(n4556), .Y(n4006) );
  OAI21X1 U3828 ( .A(n10708), .B(n10810), .C(n4449), .Y(n4007) );
  OAI21X1 U3830 ( .A(n10708), .B(n10809), .C(n6185), .Y(n4008) );
  OAI21X1 U3832 ( .A(n10708), .B(n10808), .C(n6053), .Y(n4009) );
  OAI21X1 U3834 ( .A(n10707), .B(n10807), .C(n5921), .Y(n4010) );
  OAI21X1 U3836 ( .A(n10707), .B(n10806), .C(n5662), .Y(n4011) );
  OAI21X1 U3838 ( .A(n10707), .B(n10805), .C(n4448), .Y(n4012) );
  OAI21X1 U3840 ( .A(n10707), .B(n10804), .C(n5095), .Y(n4013) );
  OAI21X1 U3842 ( .A(n10707), .B(n10803), .C(n4986), .Y(n4014) );
  OAI21X1 U3844 ( .A(n10708), .B(n10802), .C(n4877), .Y(n4015) );
  OAI21X1 U3846 ( .A(n10708), .B(n10801), .C(n4769), .Y(n4016) );
  OAI21X1 U3848 ( .A(n10708), .B(n10800), .C(n4662), .Y(n4017) );
  OAI21X1 U3850 ( .A(n10707), .B(n10799), .C(n4555), .Y(n4018) );
  OAI21X1 U3852 ( .A(n10707), .B(n10798), .C(n5203), .Y(n4019) );
  OAI21X1 U3854 ( .A(n10707), .B(n10797), .C(n6184), .Y(n4020) );
  OAI21X1 U3856 ( .A(n10707), .B(n10796), .C(n6052), .Y(n4021) );
  OAI21X1 U3858 ( .A(n10708), .B(n10795), .C(n5920), .Y(n4022) );
  OAI21X1 U3860 ( .A(n10707), .B(n10794), .C(n5789), .Y(n4023) );
  OAI21X1 U3862 ( .A(n10707), .B(n10793), .C(n5094), .Y(n4024) );
  OAI21X1 U3864 ( .A(n10707), .B(n10792), .C(n4661), .Y(n4025) );
  OAI21X1 U3866 ( .A(n10707), .B(n10791), .C(n4985), .Y(n4026) );
  OAI21X1 U3868 ( .A(n10707), .B(n10790), .C(n4876), .Y(n4027) );
  OAI21X1 U3870 ( .A(n10708), .B(n10789), .C(n4768), .Y(n4028) );
  OAI21X1 U3872 ( .A(n10708), .B(n10788), .C(n5788), .Y(n4029) );
  OAI21X1 U3874 ( .A(n10707), .B(n10787), .C(n4554), .Y(n4030) );
  OAI21X1 U3876 ( .A(n10708), .B(n10786), .C(n6183), .Y(n4031) );
  OAI21X1 U3878 ( .A(n10708), .B(n10785), .C(n5202), .Y(n4032) );
  OAI21X1 U3880 ( .A(n10707), .B(n10784), .C(n5661), .Y(n4033) );
  OAI21X1 U3882 ( .A(n10708), .B(n10783), .C(n4447), .Y(n4034) );
  OAI21X1 U3884 ( .A(n10707), .B(n10782), .C(n5544), .Y(n4035) );
  OAI21X1 U3886 ( .A(n10708), .B(n10781), .C(n5426), .Y(n4036) );
  OAI21X1 U3888 ( .A(n10708), .B(n10780), .C(n5308), .Y(n4037) );
  OAI21X1 U3890 ( .A(n10708), .B(n10779), .C(n4266), .Y(n4038) );
  OAI21X1 U3892 ( .A(n10707), .B(n10778), .C(n4265), .Y(n4039) );
  OAI21X1 U3894 ( .A(n10707), .B(n10777), .C(n5425), .Y(n4040) );
  OAI21X1 U3896 ( .A(n10707), .B(n10776), .C(n4264), .Y(n4041) );
  OAI21X1 U3898 ( .A(n10708), .B(n10775), .C(n4263), .Y(n4042) );
  OAI21X1 U3900 ( .A(n10708), .B(n10774), .C(n5919), .Y(n4043) );
  OAI21X1 U3902 ( .A(n10707), .B(n10773), .C(n5660), .Y(n4044) );
  OAI21X1 U3904 ( .A(n10708), .B(n10772), .C(n5543), .Y(n4045) );
  OAI21X1 U3906 ( .A(n10707), .B(n10771), .C(n5787), .Y(n4046) );
  OAI21X1 U3908 ( .A(n10707), .B(n10770), .C(n4262), .Y(n4047) );
  OAI21X1 U3910 ( .A(n10707), .B(n10769), .C(n5424), .Y(n4048) );
  OAI21X1 U3912 ( .A(n10708), .B(n10768), .C(n4261), .Y(n4049) );
  OAI21X1 U3914 ( .A(n10708), .B(n10767), .C(n6051), .Y(n4050) );
  OAI21X1 U3916 ( .A(n5771), .B(n6038), .C(reset_n), .Y(n1999) );
  NAND3X1 U3917 ( .A(waddr[0]), .B(n10833), .C(waddr[1]), .Y(n432) );
  OAI21X1 U3918 ( .A(n10705), .B(n10830), .C(n5093), .Y(n4051) );
  OAI21X1 U3920 ( .A(n10705), .B(n10829), .C(n5092), .Y(n4052) );
  OAI21X1 U3922 ( .A(n10705), .B(n10828), .C(n5201), .Y(n4053) );
  OAI21X1 U3924 ( .A(n10705), .B(n10827), .C(n4875), .Y(n4054) );
  OAI21X1 U3926 ( .A(n10705), .B(n10826), .C(n4984), .Y(n4055) );
  OAI21X1 U3928 ( .A(n10705), .B(n10825), .C(n4660), .Y(n4056) );
  OAI21X1 U3930 ( .A(n10705), .B(n10824), .C(n4767), .Y(n4057) );
  OAI21X1 U3932 ( .A(n10705), .B(n10823), .C(n4446), .Y(n4058) );
  OAI21X1 U3934 ( .A(n10705), .B(n10822), .C(n4553), .Y(n4059) );
  OAI21X1 U3936 ( .A(n10705), .B(n10821), .C(n6050), .Y(n4060) );
  OAI21X1 U3938 ( .A(n10705), .B(n10820), .C(n6182), .Y(n4061) );
  OAI21X1 U3940 ( .A(n10705), .B(n10819), .C(n5786), .Y(n4062) );
  OAI21X1 U3942 ( .A(n10705), .B(n10818), .C(n5918), .Y(n4063) );
  OAI21X1 U3944 ( .A(n10705), .B(n10817), .C(n5091), .Y(n4064) );
  OAI21X1 U3946 ( .A(n10705), .B(n10816), .C(n5200), .Y(n4065) );
  OAI21X1 U3948 ( .A(n10705), .B(n10815), .C(n4874), .Y(n4066) );
  OAI21X1 U3950 ( .A(n10706), .B(n10814), .C(n4983), .Y(n4067) );
  OAI21X1 U3952 ( .A(n10706), .B(n10813), .C(n4659), .Y(n4068) );
  OAI21X1 U3954 ( .A(n10705), .B(n10812), .C(n4766), .Y(n4069) );
  OAI21X1 U3956 ( .A(n10706), .B(n10811), .C(n4445), .Y(n4070) );
  OAI21X1 U3958 ( .A(n10706), .B(n10810), .C(n4552), .Y(n4071) );
  OAI21X1 U3960 ( .A(n10706), .B(n10809), .C(n6049), .Y(n4072) );
  OAI21X1 U3962 ( .A(n10706), .B(n10808), .C(n6181), .Y(n4073) );
  OAI21X1 U3964 ( .A(n10705), .B(n10807), .C(n5785), .Y(n4074) );
  OAI21X1 U3966 ( .A(n10705), .B(n10806), .C(n5542), .Y(n4075) );
  OAI21X1 U3968 ( .A(n10705), .B(n10805), .C(n4551), .Y(n4076) );
  OAI21X1 U3970 ( .A(n10705), .B(n10804), .C(n5199), .Y(n4077) );
  OAI21X1 U3972 ( .A(n10705), .B(n10803), .C(n4873), .Y(n4078) );
  OAI21X1 U3974 ( .A(n10706), .B(n10802), .C(n4982), .Y(n4079) );
  OAI21X1 U3976 ( .A(n10705), .B(n10801), .C(n4658), .Y(n4080) );
  OAI21X1 U3978 ( .A(n10706), .B(n10800), .C(n4765), .Y(n4081) );
  OAI21X1 U3980 ( .A(n10705), .B(n10799), .C(n4444), .Y(n4082) );
  OAI21X1 U3982 ( .A(n10705), .B(n10798), .C(n5090), .Y(n4083) );
  OAI21X1 U3984 ( .A(n10705), .B(n10797), .C(n6048), .Y(n4084) );
  OAI21X1 U3986 ( .A(n10706), .B(n10796), .C(n6180), .Y(n4085) );
  OAI21X1 U3988 ( .A(n10705), .B(n10795), .C(n5784), .Y(n4086) );
  OAI21X1 U3990 ( .A(n10705), .B(n10794), .C(n5917), .Y(n4087) );
  OAI21X1 U3992 ( .A(n10706), .B(n10793), .C(n5198), .Y(n4088) );
  OAI21X1 U3994 ( .A(n10705), .B(n10792), .C(n4764), .Y(n4089) );
  OAI21X1 U3996 ( .A(n10705), .B(n10791), .C(n4872), .Y(n4090) );
  OAI21X1 U3998 ( .A(n10705), .B(n10790), .C(n4981), .Y(n4091) );
  OAI21X1 U4000 ( .A(n10706), .B(n10789), .C(n4657), .Y(n4092) );
  OAI21X1 U4002 ( .A(n10706), .B(n10788), .C(n5916), .Y(n4093) );
  OAI21X1 U4004 ( .A(n10705), .B(n10787), .C(n4443), .Y(n4094) );
  OAI21X1 U4006 ( .A(n10706), .B(n10786), .C(n6047), .Y(n4095) );
  OAI21X1 U4008 ( .A(n10706), .B(n10785), .C(n5089), .Y(n4096) );
  OAI21X1 U4010 ( .A(n10705), .B(n10784), .C(n5541), .Y(n4097) );
  OAI21X1 U4012 ( .A(n10705), .B(n10783), .C(n4550), .Y(n4098) );
  OAI21X1 U4014 ( .A(n10705), .B(n10782), .C(n5659), .Y(n4099) );
  OAI21X1 U4016 ( .A(n10706), .B(n10781), .C(n5307), .Y(n4100) );
  OAI21X1 U4018 ( .A(n10706), .B(n10780), .C(n5423), .Y(n4101) );
  OAI21X1 U4020 ( .A(n10705), .B(n10779), .C(n4260), .Y(n4102) );
  OAI21X1 U4022 ( .A(n10706), .B(n10778), .C(n4259), .Y(n4103) );
  OAI21X1 U4024 ( .A(n10706), .B(n10777), .C(n5306), .Y(n4104) );
  OAI21X1 U4026 ( .A(n10705), .B(n10776), .C(n4258), .Y(n4105) );
  OAI21X1 U4028 ( .A(n10706), .B(n10775), .C(n4257), .Y(n4106) );
  OAI21X1 U4030 ( .A(n10706), .B(n10774), .C(n5783), .Y(n4107) );
  OAI21X1 U4032 ( .A(n10705), .B(n10773), .C(n5540), .Y(n4108) );
  OAI21X1 U4034 ( .A(n10706), .B(n10772), .C(n5658), .Y(n4109) );
  OAI21X1 U4036 ( .A(n10705), .B(n10771), .C(n5915), .Y(n4110) );
  OAI21X1 U4038 ( .A(n10705), .B(n10770), .C(n4256), .Y(n4111) );
  OAI21X1 U4040 ( .A(n10705), .B(n10769), .C(n5305), .Y(n4112) );
  OAI21X1 U4042 ( .A(n10706), .B(n10768), .C(n4255), .Y(n4113) );
  OAI21X1 U4044 ( .A(n10706), .B(n10767), .C(n6179), .Y(n4114) );
  OAI21X1 U4046 ( .A(n5535), .B(n6038), .C(reset_n), .Y(n2064) );
  NAND3X1 U4047 ( .A(n10835), .B(n10833), .C(waddr[1]), .Y(n498) );
  OAI21X1 U4048 ( .A(n10703), .B(n10830), .C(n4980), .Y(n4115) );
  OAI21X1 U4050 ( .A(n10703), .B(n10829), .C(n4979), .Y(n4116) );
  OAI21X1 U4052 ( .A(n10703), .B(n10828), .C(n4871), .Y(n4117) );
  OAI21X1 U4054 ( .A(n10703), .B(n10827), .C(n5197), .Y(n4118) );
  OAI21X1 U4056 ( .A(n10703), .B(n10826), .C(n5088), .Y(n4119) );
  OAI21X1 U4058 ( .A(n10703), .B(n10825), .C(n4549), .Y(n4120) );
  OAI21X1 U4060 ( .A(n10703), .B(n10824), .C(n4442), .Y(n4121) );
  OAI21X1 U4062 ( .A(n10703), .B(n10823), .C(n4763), .Y(n4122) );
  OAI21X1 U4064 ( .A(n10703), .B(n10822), .C(n4656), .Y(n4123) );
  OAI21X1 U4066 ( .A(n10703), .B(n10821), .C(n5914), .Y(n4124) );
  OAI21X1 U4068 ( .A(n10703), .B(n10820), .C(n5782), .Y(n4125) );
  OAI21X1 U4070 ( .A(n10703), .B(n10819), .C(n6178), .Y(n4126) );
  OAI21X1 U4072 ( .A(n10703), .B(n10818), .C(n6046), .Y(n4127) );
  OAI21X1 U4074 ( .A(n10703), .B(n10817), .C(n4978), .Y(n4128) );
  OAI21X1 U4076 ( .A(n10703), .B(n10816), .C(n4870), .Y(n4129) );
  OAI21X1 U4078 ( .A(n10704), .B(n10815), .C(n5196), .Y(n4130) );
  OAI21X1 U4080 ( .A(n10703), .B(n10814), .C(n5087), .Y(n4131) );
  OAI21X1 U4082 ( .A(n10704), .B(n10813), .C(n4548), .Y(n4132) );
  OAI21X1 U4084 ( .A(n10703), .B(n10812), .C(n4441), .Y(n4133) );
  OAI21X1 U4086 ( .A(n10704), .B(n10811), .C(n4762), .Y(n4134) );
  OAI21X1 U4088 ( .A(n10704), .B(n10810), .C(n4655), .Y(n4135) );
  OAI21X1 U4090 ( .A(n10704), .B(n10809), .C(n5913), .Y(n4136) );
  OAI21X1 U4092 ( .A(n10704), .B(n10808), .C(n5781), .Y(n4137) );
  OAI21X1 U4094 ( .A(n10703), .B(n10807), .C(n6177), .Y(n4138) );
  OAI21X1 U4096 ( .A(n10703), .B(n10806), .C(n5422), .Y(n4139) );
  OAI21X1 U4098 ( .A(n10703), .B(n10805), .C(n4654), .Y(n4140) );
  OAI21X1 U4100 ( .A(n10703), .B(n10804), .C(n4869), .Y(n4141) );
  OAI21X1 U4102 ( .A(n10703), .B(n10803), .C(n5195), .Y(n4142) );
  OAI21X1 U4104 ( .A(n10704), .B(n10802), .C(n5086), .Y(n4143) );
  OAI21X1 U4106 ( .A(n10704), .B(n10801), .C(n4547), .Y(n4144) );
  OAI21X1 U4108 ( .A(n10704), .B(n10800), .C(n4440), .Y(n4145) );
  OAI21X1 U4110 ( .A(n10703), .B(n10799), .C(n4761), .Y(n4146) );
  OAI21X1 U4112 ( .A(n10703), .B(n10798), .C(n4977), .Y(n4147) );
  OAI21X1 U4114 ( .A(n10703), .B(n10797), .C(n5912), .Y(n4148) );
  OAI21X1 U4116 ( .A(n10703), .B(n10796), .C(n5780), .Y(n4149) );
  OAI21X1 U4118 ( .A(n10704), .B(n10795), .C(n6176), .Y(n4150) );
  OAI21X1 U4120 ( .A(n10703), .B(n10794), .C(n6045), .Y(n4151) );
  OAI21X1 U4122 ( .A(n10703), .B(n10793), .C(n4868), .Y(n4152) );
  OAI21X1 U4124 ( .A(n10703), .B(n10792), .C(n4439), .Y(n4153) );
  OAI21X1 U4126 ( .A(n10703), .B(n10791), .C(n5194), .Y(n4154) );
  OAI21X1 U4128 ( .A(n10703), .B(n10790), .C(n5085), .Y(n4155) );
  OAI21X1 U4130 ( .A(n10704), .B(n10789), .C(n4546), .Y(n4156) );
  OAI21X1 U4132 ( .A(n10704), .B(n10788), .C(n6044), .Y(n4157) );
  OAI21X1 U4134 ( .A(n10703), .B(n10787), .C(n4760), .Y(n4158) );
  OAI21X1 U4136 ( .A(n10704), .B(n10786), .C(n5911), .Y(n4159) );
  OAI21X1 U4138 ( .A(n10704), .B(n10785), .C(n4976), .Y(n4160) );
  OAI21X1 U4140 ( .A(n10703), .B(n10784), .C(n5421), .Y(n4161) );
  OAI21X1 U4142 ( .A(n10704), .B(n10783), .C(n4653), .Y(n4162) );
  OAI21X1 U4144 ( .A(n10703), .B(n10782), .C(n5304), .Y(n4163) );
  OAI21X1 U4146 ( .A(n10704), .B(n10781), .C(n5657), .Y(n4164) );
  OAI21X1 U4148 ( .A(n10704), .B(n10780), .C(n5539), .Y(n4165) );
  OAI21X1 U4150 ( .A(n10704), .B(n10779), .C(n4254), .Y(n4166) );
  OAI21X1 U4152 ( .A(n10703), .B(n10778), .C(n4253), .Y(n4167) );
  OAI21X1 U4154 ( .A(n10703), .B(n10777), .C(n5656), .Y(n4168) );
  OAI21X1 U4156 ( .A(n10703), .B(n10776), .C(n4252), .Y(n4169) );
  OAI21X1 U4158 ( .A(n10704), .B(n10775), .C(n4251), .Y(n4170) );
  OAI21X1 U4160 ( .A(n10704), .B(n10774), .C(n6175), .Y(n4171) );
  OAI21X1 U4162 ( .A(n10703), .B(n10773), .C(n5420), .Y(n4172) );
  OAI21X1 U4164 ( .A(n10704), .B(n10772), .C(n5303), .Y(n4173) );
  OAI21X1 U4166 ( .A(n10703), .B(n10771), .C(n6043), .Y(n4174) );
  OAI21X1 U4168 ( .A(n10703), .B(n10770), .C(n4250), .Y(n4175) );
  OAI21X1 U4170 ( .A(n10703), .B(n10769), .C(n5655), .Y(n4176) );
  OAI21X1 U4172 ( .A(n10704), .B(n10768), .C(n4249), .Y(n4177) );
  OAI21X1 U4174 ( .A(n10704), .B(n10767), .C(n5779), .Y(n4178) );
  OAI21X1 U4176 ( .A(n5417), .B(n6038), .C(reset_n), .Y(n2129) );
  NAND3X1 U4177 ( .A(n10834), .B(n10833), .C(waddr[0]), .Y(n564) );
  OAI21X1 U4178 ( .A(n10701), .B(n10830), .C(n4867), .Y(n4179) );
  OAI21X1 U4181 ( .A(n10701), .B(n10829), .C(n4866), .Y(n4180) );
  OAI21X1 U4184 ( .A(n10701), .B(n10828), .C(n4975), .Y(n4181) );
  OAI21X1 U4187 ( .A(n10701), .B(n10827), .C(n5084), .Y(n4182) );
  OAI21X1 U4190 ( .A(n10701), .B(n10826), .C(n5193), .Y(n4183) );
  OAI21X1 U4193 ( .A(n10701), .B(n10825), .C(n4438), .Y(n4184) );
  OAI21X1 U4196 ( .A(n10701), .B(n10824), .C(n4545), .Y(n4185) );
  OAI21X1 U4199 ( .A(n10701), .B(n10823), .C(n4652), .Y(n4186) );
  OAI21X1 U4202 ( .A(n10701), .B(n10822), .C(n4759), .Y(n4187) );
  OAI21X1 U4205 ( .A(n10701), .B(n10821), .C(n5778), .Y(n4188) );
  OAI21X1 U4208 ( .A(n10701), .B(n10820), .C(n5910), .Y(n4189) );
  OAI21X1 U4211 ( .A(n10701), .B(n10819), .C(n6042), .Y(n4190) );
  OAI21X1 U4214 ( .A(n10701), .B(n10818), .C(n6174), .Y(n4191) );
  OAI21X1 U4217 ( .A(n10701), .B(n10817), .C(n4865), .Y(n4192) );
  OAI21X1 U4220 ( .A(n10701), .B(n10816), .C(n4974), .Y(n4193) );
  OAI21X1 U4223 ( .A(n10702), .B(n10815), .C(n5083), .Y(n4194) );
  OAI21X1 U4226 ( .A(n10701), .B(n10814), .C(n5192), .Y(n4195) );
  OAI21X1 U4229 ( .A(n10702), .B(n10813), .C(n4437), .Y(n4196) );
  OAI21X1 U4232 ( .A(n10701), .B(n10812), .C(n4544), .Y(n4197) );
  OAI21X1 U4235 ( .A(n10702), .B(n10811), .C(n4651), .Y(n4198) );
  OAI21X1 U4238 ( .A(n10702), .B(n10810), .C(n4758), .Y(n4199) );
  OAI21X1 U4241 ( .A(n10702), .B(n10809), .C(n5777), .Y(n4200) );
  OAI21X1 U4244 ( .A(n10702), .B(n10808), .C(n5909), .Y(n4201) );
  OAI21X1 U4247 ( .A(n10701), .B(n10807), .C(n6041), .Y(n4202) );
  OAI21X1 U4250 ( .A(n10701), .B(n10806), .C(n5302), .Y(n4203) );
  OAI21X1 U4253 ( .A(n10701), .B(n10805), .C(n4757), .Y(n4204) );
  OAI21X1 U4256 ( .A(n10701), .B(n10804), .C(n4973), .Y(n4205) );
  OAI21X1 U4259 ( .A(n10701), .B(n10803), .C(n5082), .Y(n4206) );
  OAI21X1 U4262 ( .A(n10702), .B(n10802), .C(n5191), .Y(n4207) );
  OAI21X1 U4265 ( .A(n10702), .B(n10801), .C(n4436), .Y(n4208) );
  OAI21X1 U4268 ( .A(n10702), .B(n10800), .C(n4543), .Y(n4209) );
  OAI21X1 U4271 ( .A(n10701), .B(n10799), .C(n4650), .Y(n4210) );
  OAI21X1 U4274 ( .A(n10701), .B(n10798), .C(n4864), .Y(n4211) );
  OAI21X1 U4277 ( .A(n10701), .B(n10797), .C(n5776), .Y(n4212) );
  OAI21X1 U4280 ( .A(n10701), .B(n10796), .C(n5908), .Y(n4213) );
  OAI21X1 U4283 ( .A(n10702), .B(n10795), .C(n6040), .Y(n4214) );
  OAI21X1 U4286 ( .A(n10701), .B(n10794), .C(n6173), .Y(n4215) );
  OAI21X1 U4289 ( .A(n10701), .B(n10793), .C(n4972), .Y(n4216) );
  OAI21X1 U4292 ( .A(n10701), .B(n10792), .C(n4542), .Y(n4217) );
  OAI21X1 U4295 ( .A(n10701), .B(n10791), .C(n5081), .Y(n4218) );
  OAI21X1 U4298 ( .A(n10701), .B(n10790), .C(n5190), .Y(n4219) );
  OAI21X1 U4301 ( .A(n10702), .B(n10789), .C(n4435), .Y(n4220) );
  OAI21X1 U4304 ( .A(n10702), .B(n10788), .C(n6172), .Y(n4221) );
  OAI21X1 U4307 ( .A(n10701), .B(n10787), .C(n4649), .Y(n4222) );
  OAI21X1 U4310 ( .A(n10702), .B(n10786), .C(n5775), .Y(n4223) );
  OAI21X1 U4313 ( .A(n10702), .B(n10785), .C(n4863), .Y(n4224) );
  OAI21X1 U4316 ( .A(n10701), .B(n10784), .C(n5301), .Y(n4225) );
  OAI21X1 U4319 ( .A(n10702), .B(n10783), .C(n4756), .Y(n4226) );
  OAI21X1 U4322 ( .A(n10701), .B(n10782), .C(n5419), .Y(n4227) );
  OAI21X1 U4325 ( .A(n10702), .B(n10781), .C(n5538), .Y(n4228) );
  OAI21X1 U4328 ( .A(n10702), .B(n10780), .C(n5654), .Y(n4229) );
  OAI21X1 U4331 ( .A(n10702), .B(n10779), .C(n4248), .Y(n4230) );
  OAI21X1 U4334 ( .A(n10701), .B(n10778), .C(n4247), .Y(n4231) );
  OAI21X1 U4337 ( .A(n10701), .B(n10777), .C(n5537), .Y(n4232) );
  OAI21X1 U4340 ( .A(n10701), .B(n10776), .C(n4246), .Y(n4233) );
  OAI21X1 U4343 ( .A(n10702), .B(n10775), .C(n4245), .Y(n4234) );
  OAI21X1 U4346 ( .A(n10702), .B(n10774), .C(n6039), .Y(n4235) );
  OAI21X1 U4349 ( .A(n10701), .B(n10773), .C(n5300), .Y(n4236) );
  OAI21X1 U4352 ( .A(n10702), .B(n10772), .C(n5418), .Y(n4237) );
  OAI21X1 U4355 ( .A(n10701), .B(n10771), .C(n6171), .Y(n4238) );
  OAI21X1 U4358 ( .A(n10701), .B(n10770), .C(n4244), .Y(n4239) );
  OAI21X1 U4361 ( .A(n10701), .B(n10769), .C(n5536), .Y(n4240) );
  OAI21X1 U4364 ( .A(n10702), .B(n10768), .C(n4243), .Y(n4241) );
  OAI21X1 U4367 ( .A(n10702), .B(n10767), .C(n5907), .Y(n4242) );
  OAI21X1 U4370 ( .A(n5299), .B(n6038), .C(reset_n), .Y(n2194) );
  NAND3X1 U4371 ( .A(n10832), .B(n10831), .C(n631), .Y(n1739) );
  NAND3X1 U4372 ( .A(n10834), .B(n10833), .C(n10835), .Y(n630) );
  AND2X1 U4373 ( .A(\RF[0][62] ), .B(n10702), .Y(n2192) );
  INVX1 U4374 ( .A(n2192), .Y(n4243) );
  AND2X1 U4375 ( .A(\RF[0][60] ), .B(n10702), .Y(n2190) );
  INVX1 U4376 ( .A(n2190), .Y(n4244) );
  AND2X1 U4377 ( .A(\RF[0][55] ), .B(n10701), .Y(n2185) );
  INVX1 U4378 ( .A(n2185), .Y(n4245) );
  AND2X1 U4379 ( .A(\RF[0][54] ), .B(n10702), .Y(n2184) );
  INVX1 U4380 ( .A(n2184), .Y(n4246) );
  AND2X1 U4381 ( .A(\RF[0][52] ), .B(n10701), .Y(n2182) );
  INVX1 U4382 ( .A(n2182), .Y(n4247) );
  AND2X1 U4383 ( .A(\RF[0][51] ), .B(n10702), .Y(n2181) );
  INVX1 U4384 ( .A(n2181), .Y(n4248) );
  AND2X1 U4385 ( .A(\RF[1][62] ), .B(n10704), .Y(n2127) );
  INVX1 U4386 ( .A(n2127), .Y(n4249) );
  AND2X1 U4387 ( .A(\RF[1][60] ), .B(n10704), .Y(n2125) );
  INVX1 U4388 ( .A(n2125), .Y(n4250) );
  AND2X1 U4389 ( .A(\RF[1][55] ), .B(n10703), .Y(n2120) );
  INVX1 U4390 ( .A(n2120), .Y(n4251) );
  AND2X1 U4391 ( .A(\RF[1][54] ), .B(n10704), .Y(n2119) );
  INVX1 U4392 ( .A(n2119), .Y(n4252) );
  AND2X1 U4393 ( .A(\RF[1][52] ), .B(n10703), .Y(n2117) );
  INVX1 U4394 ( .A(n2117), .Y(n4253) );
  AND2X1 U4395 ( .A(\RF[1][51] ), .B(n10704), .Y(n2116) );
  INVX1 U4396 ( .A(n2116), .Y(n4254) );
  AND2X1 U4397 ( .A(\RF[2][62] ), .B(n10706), .Y(n2062) );
  INVX1 U4398 ( .A(n2062), .Y(n4255) );
  AND2X1 U4399 ( .A(\RF[2][60] ), .B(n10705), .Y(n2060) );
  INVX1 U4400 ( .A(n2060), .Y(n4256) );
  AND2X1 U4401 ( .A(\RF[2][55] ), .B(n10705), .Y(n2055) );
  INVX1 U4402 ( .A(n2055), .Y(n4257) );
  AND2X1 U4403 ( .A(\RF[2][54] ), .B(n10706), .Y(n2054) );
  INVX1 U4404 ( .A(n2054), .Y(n4258) );
  AND2X1 U4405 ( .A(\RF[2][52] ), .B(n10706), .Y(n2052) );
  INVX1 U4406 ( .A(n2052), .Y(n4259) );
  AND2X1 U4407 ( .A(\RF[2][51] ), .B(n10706), .Y(n2051) );
  INVX1 U4408 ( .A(n2051), .Y(n4260) );
  AND2X1 U4409 ( .A(\RF[3][62] ), .B(n10707), .Y(n1997) );
  INVX1 U4410 ( .A(n1997), .Y(n4261) );
  AND2X1 U4411 ( .A(\RF[3][60] ), .B(n10708), .Y(n1995) );
  INVX1 U4412 ( .A(n1995), .Y(n4262) );
  AND2X1 U4413 ( .A(\RF[3][55] ), .B(n10708), .Y(n1990) );
  INVX1 U4414 ( .A(n1990), .Y(n4263) );
  AND2X1 U4415 ( .A(\RF[3][54] ), .B(n10708), .Y(n1989) );
  INVX1 U4416 ( .A(n1989), .Y(n4264) );
  AND2X1 U4417 ( .A(\RF[3][52] ), .B(n10707), .Y(n1987) );
  INVX1 U4418 ( .A(n1987), .Y(n4265) );
  AND2X1 U4419 ( .A(\RF[3][51] ), .B(n10708), .Y(n1986) );
  INVX1 U4420 ( .A(n1986), .Y(n4266) );
  AND2X1 U4421 ( .A(\RF[4][62] ), .B(n10709), .Y(n1932) );
  INVX1 U4422 ( .A(n1932), .Y(n4267) );
  AND2X1 U4423 ( .A(\RF[4][60] ), .B(n10710), .Y(n1930) );
  INVX1 U4424 ( .A(n1930), .Y(n4268) );
  AND2X1 U4425 ( .A(\RF[4][55] ), .B(n10710), .Y(n1925) );
  INVX1 U4426 ( .A(n1925), .Y(n4269) );
  AND2X1 U4427 ( .A(\RF[4][54] ), .B(n10710), .Y(n1924) );
  INVX1 U4428 ( .A(n1924), .Y(n4270) );
  AND2X1 U4429 ( .A(\RF[4][52] ), .B(n10709), .Y(n1922) );
  INVX1 U4430 ( .A(n1922), .Y(n4271) );
  AND2X1 U4431 ( .A(\RF[4][51] ), .B(n10710), .Y(n1921) );
  INVX1 U4432 ( .A(n1921), .Y(n4272) );
  AND2X1 U4433 ( .A(\RF[5][62] ), .B(n10712), .Y(n1867) );
  INVX1 U4434 ( .A(n1867), .Y(n4273) );
  AND2X1 U4435 ( .A(\RF[5][60] ), .B(n10711), .Y(n1865) );
  INVX1 U4436 ( .A(n1865), .Y(n4274) );
  AND2X1 U4437 ( .A(\RF[5][55] ), .B(n10711), .Y(n1860) );
  INVX1 U4438 ( .A(n1860), .Y(n4275) );
  AND2X1 U4439 ( .A(\RF[5][54] ), .B(n10712), .Y(n1859) );
  INVX1 U4440 ( .A(n1859), .Y(n4276) );
  AND2X1 U4441 ( .A(\RF[5][52] ), .B(n10712), .Y(n1857) );
  INVX1 U4442 ( .A(n1857), .Y(n4277) );
  AND2X1 U4443 ( .A(\RF[5][51] ), .B(n10712), .Y(n1856) );
  INVX1 U4444 ( .A(n1856), .Y(n4278) );
  AND2X1 U4445 ( .A(\RF[6][62] ), .B(n10714), .Y(n1802) );
  INVX1 U4446 ( .A(n1802), .Y(n4279) );
  AND2X1 U4447 ( .A(\RF[6][60] ), .B(n10713), .Y(n1800) );
  INVX1 U4448 ( .A(n1800), .Y(n4280) );
  AND2X1 U4449 ( .A(\RF[6][55] ), .B(n10713), .Y(n1795) );
  INVX1 U4450 ( .A(n1795), .Y(n4281) );
  AND2X1 U4451 ( .A(\RF[6][54] ), .B(n10714), .Y(n1794) );
  INVX1 U4452 ( .A(n1794), .Y(n4282) );
  AND2X1 U4453 ( .A(\RF[6][52] ), .B(n10714), .Y(n1792) );
  INVX1 U4454 ( .A(n1792), .Y(n4283) );
  AND2X1 U4455 ( .A(\RF[6][51] ), .B(n10714), .Y(n1791) );
  INVX1 U4456 ( .A(n1791), .Y(n4284) );
  AND2X1 U4457 ( .A(\RF[7][62] ), .B(n10716), .Y(n1736) );
  INVX1 U4458 ( .A(n1736), .Y(n4285) );
  AND2X1 U4459 ( .A(\RF[7][60] ), .B(n10715), .Y(n1734) );
  INVX1 U4460 ( .A(n1734), .Y(n4286) );
  AND2X1 U4461 ( .A(\RF[7][55] ), .B(n10715), .Y(n1729) );
  INVX1 U4462 ( .A(n1729), .Y(n4287) );
  AND2X1 U4463 ( .A(\RF[7][54] ), .B(n10716), .Y(n1728) );
  INVX1 U4464 ( .A(n1728), .Y(n4288) );
  AND2X1 U4465 ( .A(\RF[7][52] ), .B(n10716), .Y(n1726) );
  INVX1 U4466 ( .A(n1726), .Y(n4289) );
  AND2X1 U4467 ( .A(\RF[7][51] ), .B(n10716), .Y(n1725) );
  INVX1 U4468 ( .A(n1725), .Y(n4290) );
  AND2X1 U4469 ( .A(\RF[8][62] ), .B(n10718), .Y(n1671) );
  INVX1 U4470 ( .A(n1671), .Y(n4291) );
  AND2X1 U4471 ( .A(\RF[8][60] ), .B(n10717), .Y(n1669) );
  INVX1 U4472 ( .A(n1669), .Y(n4292) );
  AND2X1 U4473 ( .A(\RF[8][55] ), .B(n10717), .Y(n1664) );
  INVX1 U4474 ( .A(n1664), .Y(n4293) );
  AND2X1 U4475 ( .A(\RF[8][54] ), .B(n10718), .Y(n1663) );
  INVX1 U4476 ( .A(n1663), .Y(n4294) );
  AND2X1 U4477 ( .A(\RF[8][52] ), .B(n10718), .Y(n1661) );
  INVX1 U4478 ( .A(n1661), .Y(n4295) );
  AND2X1 U4479 ( .A(\RF[8][51] ), .B(n10718), .Y(n1660) );
  INVX1 U4480 ( .A(n1660), .Y(n4296) );
  AND2X1 U4481 ( .A(\RF[9][62] ), .B(n10720), .Y(n1606) );
  INVX1 U4482 ( .A(n1606), .Y(n4297) );
  AND2X1 U4483 ( .A(\RF[9][60] ), .B(n10719), .Y(n1604) );
  INVX1 U4484 ( .A(n1604), .Y(n4298) );
  AND2X1 U4485 ( .A(\RF[9][55] ), .B(n10719), .Y(n1599) );
  INVX1 U4486 ( .A(n1599), .Y(n4299) );
  AND2X1 U4487 ( .A(\RF[9][54] ), .B(n10720), .Y(n1598) );
  INVX1 U4488 ( .A(n1598), .Y(n4300) );
  AND2X1 U4489 ( .A(\RF[9][52] ), .B(n10720), .Y(n1596) );
  INVX1 U4490 ( .A(n1596), .Y(n4301) );
  AND2X1 U4491 ( .A(\RF[9][51] ), .B(n10720), .Y(n1595) );
  INVX1 U4492 ( .A(n1595), .Y(n4302) );
  AND2X1 U4493 ( .A(\RF[10][62] ), .B(n10722), .Y(n1541) );
  INVX1 U4494 ( .A(n1541), .Y(n4303) );
  AND2X1 U4495 ( .A(\RF[10][60] ), .B(n10721), .Y(n1539) );
  INVX1 U4496 ( .A(n1539), .Y(n4304) );
  AND2X1 U4497 ( .A(\RF[10][55] ), .B(n10721), .Y(n1534) );
  INVX1 U4498 ( .A(n1534), .Y(n4305) );
  AND2X1 U4499 ( .A(\RF[10][54] ), .B(n10722), .Y(n1533) );
  INVX1 U4500 ( .A(n1533), .Y(n4306) );
  AND2X1 U4501 ( .A(\RF[10][52] ), .B(n10722), .Y(n1531) );
  INVX1 U4502 ( .A(n1531), .Y(n4307) );
  AND2X1 U4503 ( .A(\RF[10][51] ), .B(n10722), .Y(n1530) );
  INVX1 U4504 ( .A(n1530), .Y(n4308) );
  AND2X1 U4505 ( .A(\RF[11][62] ), .B(n10724), .Y(n1476) );
  INVX1 U4506 ( .A(n1476), .Y(n4309) );
  AND2X1 U4507 ( .A(\RF[11][60] ), .B(n10723), .Y(n1474) );
  INVX1 U4508 ( .A(n1474), .Y(n4310) );
  AND2X1 U4509 ( .A(\RF[11][55] ), .B(n10723), .Y(n1469) );
  INVX1 U4510 ( .A(n1469), .Y(n4311) );
  AND2X1 U4511 ( .A(\RF[11][54] ), .B(n10724), .Y(n1468) );
  INVX1 U4512 ( .A(n1468), .Y(n4312) );
  AND2X1 U4513 ( .A(\RF[11][52] ), .B(n10724), .Y(n1466) );
  INVX1 U4514 ( .A(n1466), .Y(n4313) );
  AND2X1 U4515 ( .A(\RF[11][51] ), .B(n10724), .Y(n1465) );
  INVX1 U4516 ( .A(n1465), .Y(n4314) );
  AND2X1 U4517 ( .A(\RF[12][62] ), .B(n10726), .Y(n1411) );
  INVX1 U4518 ( .A(n1411), .Y(n4315) );
  AND2X1 U4519 ( .A(\RF[12][60] ), .B(n10726), .Y(n1409) );
  INVX1 U4520 ( .A(n1409), .Y(n4316) );
  AND2X1 U4521 ( .A(\RF[12][55] ), .B(n10725), .Y(n1404) );
  INVX1 U4522 ( .A(n1404), .Y(n4317) );
  AND2X1 U4523 ( .A(\RF[12][54] ), .B(n10726), .Y(n1403) );
  INVX1 U4524 ( .A(n1403), .Y(n4318) );
  AND2X1 U4525 ( .A(\RF[12][52] ), .B(n10725), .Y(n1401) );
  INVX1 U4526 ( .A(n1401), .Y(n4319) );
  AND2X1 U4527 ( .A(\RF[12][51] ), .B(n10726), .Y(n1400) );
  INVX1 U4528 ( .A(n1400), .Y(n4320) );
  AND2X1 U4529 ( .A(\RF[13][62] ), .B(n10728), .Y(n1346) );
  INVX1 U4530 ( .A(n1346), .Y(n4321) );
  AND2X1 U4531 ( .A(\RF[13][60] ), .B(n10728), .Y(n1344) );
  INVX1 U4532 ( .A(n1344), .Y(n4322) );
  AND2X1 U4533 ( .A(\RF[13][55] ), .B(n10727), .Y(n1339) );
  INVX1 U4534 ( .A(n1339), .Y(n4323) );
  AND2X1 U4535 ( .A(\RF[13][54] ), .B(n10728), .Y(n1338) );
  INVX1 U4536 ( .A(n1338), .Y(n4324) );
  AND2X1 U4537 ( .A(\RF[13][52] ), .B(n10727), .Y(n1336) );
  INVX1 U4538 ( .A(n1336), .Y(n4325) );
  AND2X1 U4539 ( .A(\RF[13][51] ), .B(n10728), .Y(n1335) );
  INVX1 U4540 ( .A(n1335), .Y(n4326) );
  AND2X1 U4541 ( .A(\RF[14][62] ), .B(n10730), .Y(n1281) );
  INVX1 U4542 ( .A(n1281), .Y(n4327) );
  AND2X1 U4543 ( .A(\RF[14][60] ), .B(n10729), .Y(n1279) );
  INVX1 U4544 ( .A(n1279), .Y(n4328) );
  AND2X1 U4545 ( .A(\RF[14][55] ), .B(n10729), .Y(n1274) );
  INVX1 U4546 ( .A(n1274), .Y(n4329) );
  AND2X1 U4547 ( .A(\RF[14][54] ), .B(n10730), .Y(n1273) );
  INVX1 U4548 ( .A(n1273), .Y(n4330) );
  AND2X1 U4549 ( .A(\RF[14][52] ), .B(n10730), .Y(n1271) );
  INVX1 U4550 ( .A(n1271), .Y(n4331) );
  AND2X1 U4551 ( .A(\RF[14][51] ), .B(n10730), .Y(n1270) );
  INVX1 U4552 ( .A(n1270), .Y(n4332) );
  AND2X1 U4553 ( .A(\RF[15][62] ), .B(n10731), .Y(n1215) );
  INVX1 U4554 ( .A(n1215), .Y(n4333) );
  AND2X1 U4555 ( .A(\RF[15][60] ), .B(n10732), .Y(n1213) );
  INVX1 U4556 ( .A(n1213), .Y(n4334) );
  AND2X1 U4557 ( .A(\RF[15][55] ), .B(n10732), .Y(n1208) );
  INVX1 U4558 ( .A(n1208), .Y(n4335) );
  AND2X1 U4559 ( .A(\RF[15][54] ), .B(n10732), .Y(n1207) );
  INVX1 U4560 ( .A(n1207), .Y(n4336) );
  AND2X1 U4561 ( .A(\RF[15][52] ), .B(n10731), .Y(n1205) );
  INVX1 U4562 ( .A(n1205), .Y(n4337) );
  AND2X1 U4563 ( .A(\RF[15][51] ), .B(n10732), .Y(n1204) );
  INVX1 U4564 ( .A(n1204), .Y(n4338) );
  AND2X1 U4565 ( .A(\RF[16][62] ), .B(n10733), .Y(n1150) );
  INVX1 U4566 ( .A(n1150), .Y(n4339) );
  AND2X1 U4567 ( .A(\RF[16][60] ), .B(n10734), .Y(n1148) );
  INVX1 U4568 ( .A(n1148), .Y(n4340) );
  AND2X1 U4569 ( .A(\RF[16][55] ), .B(n10734), .Y(n1143) );
  INVX1 U4570 ( .A(n1143), .Y(n4341) );
  AND2X1 U4571 ( .A(\RF[16][54] ), .B(n10734), .Y(n1142) );
  INVX1 U4572 ( .A(n1142), .Y(n4342) );
  AND2X1 U4573 ( .A(\RF[16][52] ), .B(n10733), .Y(n1140) );
  INVX1 U4574 ( .A(n1140), .Y(n4343) );
  AND2X1 U4575 ( .A(\RF[16][51] ), .B(n10734), .Y(n1139) );
  INVX1 U4576 ( .A(n1139), .Y(n4344) );
  AND2X1 U4577 ( .A(\RF[17][62] ), .B(n10736), .Y(n1085) );
  INVX1 U4578 ( .A(n1085), .Y(n4345) );
  AND2X1 U4579 ( .A(\RF[17][60] ), .B(n10735), .Y(n1083) );
  INVX1 U4580 ( .A(n1083), .Y(n4346) );
  AND2X1 U4581 ( .A(\RF[17][55] ), .B(n10735), .Y(n1078) );
  INVX1 U4582 ( .A(n1078), .Y(n4347) );
  AND2X1 U4583 ( .A(\RF[17][54] ), .B(n10736), .Y(n1077) );
  INVX1 U4584 ( .A(n1077), .Y(n4348) );
  AND2X1 U4585 ( .A(\RF[17][52] ), .B(n10736), .Y(n1075) );
  INVX1 U4586 ( .A(n1075), .Y(n4349) );
  AND2X1 U4587 ( .A(\RF[17][51] ), .B(n10736), .Y(n1074) );
  INVX1 U4588 ( .A(n1074), .Y(n4350) );
  AND2X1 U4589 ( .A(\RF[18][62] ), .B(n10738), .Y(n1020) );
  INVX1 U4590 ( .A(n1020), .Y(n4351) );
  AND2X1 U4591 ( .A(\RF[18][60] ), .B(n10737), .Y(n1018) );
  INVX1 U4592 ( .A(n1018), .Y(n4352) );
  AND2X1 U4593 ( .A(\RF[18][55] ), .B(n10737), .Y(n1013) );
  INVX1 U4594 ( .A(n1013), .Y(n4353) );
  AND2X1 U4595 ( .A(\RF[18][54] ), .B(n10738), .Y(n1012) );
  INVX1 U4596 ( .A(n1012), .Y(n4354) );
  AND2X1 U4597 ( .A(\RF[18][52] ), .B(n10738), .Y(n1010) );
  INVX1 U4598 ( .A(n1010), .Y(n4355) );
  AND2X1 U4599 ( .A(\RF[18][51] ), .B(n10738), .Y(n1009) );
  INVX1 U4600 ( .A(n1009), .Y(n4356) );
  AND2X1 U4601 ( .A(\RF[19][62] ), .B(n10740), .Y(n955) );
  INVX1 U4602 ( .A(n955), .Y(n4357) );
  AND2X1 U4603 ( .A(\RF[19][60] ), .B(n10739), .Y(n953) );
  INVX1 U4604 ( .A(n953), .Y(n4358) );
  AND2X1 U4605 ( .A(\RF[19][55] ), .B(n10739), .Y(n948) );
  INVX1 U4606 ( .A(n948), .Y(n4359) );
  AND2X1 U4607 ( .A(\RF[19][54] ), .B(n10740), .Y(n947) );
  INVX1 U4608 ( .A(n947), .Y(n4360) );
  AND2X1 U4609 ( .A(\RF[19][52] ), .B(n10740), .Y(n945) );
  INVX1 U4610 ( .A(n945), .Y(n4361) );
  AND2X1 U4611 ( .A(\RF[19][51] ), .B(n10740), .Y(n944) );
  INVX1 U4612 ( .A(n944), .Y(n4362) );
  AND2X1 U4613 ( .A(\RF[20][62] ), .B(n10742), .Y(n890) );
  INVX1 U4614 ( .A(n890), .Y(n4363) );
  AND2X1 U4615 ( .A(\RF[20][60] ), .B(n10741), .Y(n888) );
  INVX1 U4616 ( .A(n888), .Y(n4364) );
  AND2X1 U4617 ( .A(\RF[20][55] ), .B(n10741), .Y(n883) );
  INVX1 U4618 ( .A(n883), .Y(n4365) );
  AND2X1 U4619 ( .A(\RF[20][54] ), .B(n10742), .Y(n882) );
  INVX1 U4620 ( .A(n882), .Y(n4366) );
  AND2X1 U4621 ( .A(\RF[20][52] ), .B(n10742), .Y(n880) );
  INVX1 U4622 ( .A(n880), .Y(n4367) );
  AND2X1 U4623 ( .A(\RF[20][51] ), .B(n10742), .Y(n879) );
  INVX1 U4624 ( .A(n879), .Y(n4368) );
  AND2X1 U4625 ( .A(\RF[21][62] ), .B(n10744), .Y(n825) );
  INVX1 U4626 ( .A(n825), .Y(n4369) );
  AND2X1 U4627 ( .A(\RF[21][60] ), .B(n10743), .Y(n823) );
  INVX1 U4628 ( .A(n823), .Y(n4370) );
  AND2X1 U4629 ( .A(\RF[21][55] ), .B(n10743), .Y(n818) );
  INVX1 U4630 ( .A(n818), .Y(n4371) );
  AND2X1 U4631 ( .A(\RF[21][54] ), .B(n10744), .Y(n817) );
  INVX1 U4632 ( .A(n817), .Y(n4372) );
  AND2X1 U4633 ( .A(\RF[21][52] ), .B(n10744), .Y(n815) );
  INVX1 U4634 ( .A(n815), .Y(n4373) );
  AND2X1 U4635 ( .A(\RF[21][51] ), .B(n10744), .Y(n814) );
  INVX1 U4636 ( .A(n814), .Y(n4374) );
  AND2X1 U4637 ( .A(\RF[22][62] ), .B(n10746), .Y(n760) );
  INVX1 U4638 ( .A(n760), .Y(n4375) );
  AND2X1 U4639 ( .A(\RF[22][60] ), .B(n10745), .Y(n758) );
  INVX1 U4640 ( .A(n758), .Y(n4376) );
  AND2X1 U4641 ( .A(\RF[22][55] ), .B(n10745), .Y(n753) );
  INVX1 U4642 ( .A(n753), .Y(n4377) );
  AND2X1 U4643 ( .A(\RF[22][54] ), .B(n10746), .Y(n752) );
  INVX1 U4644 ( .A(n752), .Y(n4378) );
  AND2X1 U4645 ( .A(\RF[22][52] ), .B(n10746), .Y(n750) );
  INVX1 U4646 ( .A(n750), .Y(n4379) );
  AND2X1 U4647 ( .A(\RF[22][51] ), .B(n10746), .Y(n749) );
  INVX1 U4648 ( .A(n749), .Y(n4380) );
  AND2X1 U4649 ( .A(\RF[23][62] ), .B(n10748), .Y(n694) );
  INVX1 U4650 ( .A(n694), .Y(n4381) );
  AND2X1 U4651 ( .A(\RF[23][60] ), .B(n10747), .Y(n692) );
  INVX1 U4652 ( .A(n692), .Y(n4382) );
  AND2X1 U4653 ( .A(\RF[23][55] ), .B(n10747), .Y(n687) );
  INVX1 U4654 ( .A(n687), .Y(n4383) );
  AND2X1 U4655 ( .A(\RF[23][54] ), .B(n10748), .Y(n686) );
  INVX1 U4656 ( .A(n686), .Y(n4384) );
  AND2X1 U4657 ( .A(\RF[23][52] ), .B(n10748), .Y(n684) );
  INVX1 U4658 ( .A(n684), .Y(n4385) );
  AND2X1 U4659 ( .A(\RF[23][51] ), .B(n10748), .Y(n683) );
  INVX1 U4660 ( .A(n683), .Y(n4386) );
  AND2X1 U4661 ( .A(\RF[24][62] ), .B(n10749), .Y(n627) );
  INVX1 U4662 ( .A(n627), .Y(n4387) );
  AND2X1 U4663 ( .A(\RF[24][60] ), .B(n10750), .Y(n625) );
  INVX1 U4664 ( .A(n625), .Y(n4388) );
  AND2X1 U4665 ( .A(\RF[24][55] ), .B(n10750), .Y(n620) );
  INVX1 U4666 ( .A(n620), .Y(n4389) );
  AND2X1 U4667 ( .A(\RF[24][54] ), .B(n10750), .Y(n619) );
  INVX1 U4668 ( .A(n619), .Y(n4390) );
  AND2X1 U4669 ( .A(\RF[24][52] ), .B(n10749), .Y(n617) );
  INVX1 U4670 ( .A(n617), .Y(n4391) );
  AND2X1 U4671 ( .A(\RF[24][51] ), .B(n10750), .Y(n616) );
  INVX1 U4672 ( .A(n616), .Y(n4392) );
  AND2X1 U4673 ( .A(\RF[25][62] ), .B(n10752), .Y(n561) );
  INVX1 U4674 ( .A(n561), .Y(n4393) );
  AND2X1 U4675 ( .A(\RF[25][60] ), .B(n10751), .Y(n559) );
  INVX1 U4676 ( .A(n559), .Y(n4394) );
  AND2X1 U4677 ( .A(\RF[25][55] ), .B(n10751), .Y(n554) );
  INVX1 U4678 ( .A(n554), .Y(n4395) );
  AND2X1 U4679 ( .A(\RF[25][54] ), .B(n10752), .Y(n553) );
  INVX1 U4680 ( .A(n553), .Y(n4396) );
  AND2X1 U4681 ( .A(\RF[25][52] ), .B(n10752), .Y(n551) );
  INVX1 U4682 ( .A(n551), .Y(n4397) );
  AND2X1 U4683 ( .A(\RF[25][51] ), .B(n10752), .Y(n550) );
  INVX1 U4684 ( .A(n550), .Y(n4398) );
  AND2X1 U4685 ( .A(\RF[26][62] ), .B(n10754), .Y(n495) );
  INVX1 U4686 ( .A(n495), .Y(n4399) );
  AND2X1 U4687 ( .A(\RF[26][60] ), .B(n10753), .Y(n493) );
  INVX1 U4688 ( .A(n493), .Y(n4400) );
  AND2X1 U4689 ( .A(\RF[26][55] ), .B(n10753), .Y(n488) );
  INVX1 U4690 ( .A(n488), .Y(n4401) );
  AND2X1 U4691 ( .A(\RF[26][54] ), .B(n10754), .Y(n487) );
  INVX1 U4692 ( .A(n487), .Y(n4402) );
  AND2X1 U4693 ( .A(\RF[26][52] ), .B(n10754), .Y(n485) );
  INVX1 U4694 ( .A(n485), .Y(n4403) );
  AND2X1 U4695 ( .A(\RF[26][51] ), .B(n10754), .Y(n484) );
  INVX1 U4696 ( .A(n484), .Y(n4404) );
  AND2X1 U4697 ( .A(\RF[27][62] ), .B(n10756), .Y(n429) );
  INVX1 U4698 ( .A(n429), .Y(n4405) );
  AND2X1 U4699 ( .A(\RF[27][60] ), .B(n10755), .Y(n427) );
  INVX1 U4700 ( .A(n427), .Y(n4406) );
  AND2X1 U4701 ( .A(\RF[27][55] ), .B(n10755), .Y(n422) );
  INVX1 U4702 ( .A(n422), .Y(n4407) );
  AND2X1 U4703 ( .A(\RF[27][54] ), .B(n10756), .Y(n421) );
  INVX1 U4704 ( .A(n421), .Y(n4408) );
  AND2X1 U4705 ( .A(\RF[27][52] ), .B(n10756), .Y(n419) );
  INVX1 U4706 ( .A(n419), .Y(n4409) );
  AND2X1 U4707 ( .A(\RF[27][51] ), .B(n10756), .Y(n418) );
  INVX1 U4708 ( .A(n418), .Y(n4410) );
  AND2X1 U4709 ( .A(\RF[28][62] ), .B(n10758), .Y(n363) );
  INVX1 U4710 ( .A(n363), .Y(n4411) );
  AND2X1 U4711 ( .A(\RF[28][60] ), .B(n10757), .Y(n361) );
  INVX1 U4712 ( .A(n361), .Y(n4412) );
  AND2X1 U4713 ( .A(\RF[28][55] ), .B(n10757), .Y(n356) );
  INVX1 U4714 ( .A(n356), .Y(n4413) );
  AND2X1 U4715 ( .A(\RF[28][54] ), .B(n10758), .Y(n355) );
  INVX1 U4716 ( .A(n355), .Y(n4414) );
  AND2X1 U4717 ( .A(\RF[28][52] ), .B(n10758), .Y(n353) );
  INVX1 U4718 ( .A(n353), .Y(n4415) );
  AND2X1 U4719 ( .A(\RF[28][51] ), .B(n10758), .Y(n352) );
  INVX1 U4720 ( .A(n352), .Y(n4416) );
  AND2X1 U4721 ( .A(\RF[29][62] ), .B(n10760), .Y(n297) );
  INVX1 U4722 ( .A(n297), .Y(n4417) );
  AND2X1 U4723 ( .A(\RF[29][60] ), .B(n10759), .Y(n295) );
  INVX1 U4724 ( .A(n295), .Y(n4418) );
  AND2X1 U4725 ( .A(\RF[29][55] ), .B(n10759), .Y(n290) );
  INVX1 U4726 ( .A(n290), .Y(n4419) );
  AND2X1 U4727 ( .A(\RF[29][54] ), .B(n10760), .Y(n289) );
  INVX1 U4728 ( .A(n289), .Y(n4420) );
  AND2X1 U4729 ( .A(\RF[29][52] ), .B(n10760), .Y(n287) );
  INVX1 U4730 ( .A(n287), .Y(n4421) );
  AND2X1 U4731 ( .A(\RF[29][51] ), .B(n10760), .Y(n286) );
  INVX1 U4732 ( .A(n286), .Y(n4422) );
  AND2X1 U4733 ( .A(\RF[30][62] ), .B(n10762), .Y(n231) );
  INVX1 U4734 ( .A(n231), .Y(n4423) );
  AND2X1 U4735 ( .A(\RF[30][60] ), .B(n10761), .Y(n229) );
  INVX1 U4736 ( .A(n229), .Y(n4424) );
  AND2X1 U4737 ( .A(\RF[30][55] ), .B(n10761), .Y(n224) );
  INVX1 U4738 ( .A(n224), .Y(n4425) );
  AND2X1 U4739 ( .A(\RF[30][54] ), .B(n10762), .Y(n223) );
  INVX1 U4740 ( .A(n223), .Y(n4426) );
  AND2X1 U4741 ( .A(\RF[30][52] ), .B(n10762), .Y(n221) );
  INVX1 U4742 ( .A(n221), .Y(n4427) );
  AND2X1 U4743 ( .A(\RF[30][51] ), .B(n10762), .Y(n220) );
  INVX1 U4744 ( .A(n220), .Y(n4428) );
  AND2X1 U4745 ( .A(\RF[31][62] ), .B(n10764), .Y(n163) );
  INVX1 U4746 ( .A(n163), .Y(n4429) );
  AND2X1 U4747 ( .A(\RF[31][60] ), .B(n10763), .Y(n159) );
  INVX1 U4748 ( .A(n159), .Y(n4430) );
  AND2X1 U4749 ( .A(\RF[31][55] ), .B(n10763), .Y(n149) );
  INVX1 U4750 ( .A(n149), .Y(n4431) );
  AND2X1 U4751 ( .A(\RF[31][54] ), .B(n10764), .Y(n147) );
  INVX1 U4752 ( .A(n147), .Y(n4432) );
  AND2X1 U4753 ( .A(\RF[31][52] ), .B(n10764), .Y(n143) );
  INVX1 U4754 ( .A(n143), .Y(n4433) );
  AND2X1 U4755 ( .A(\RF[31][51] ), .B(n10764), .Y(n141) );
  INVX1 U4756 ( .A(n141), .Y(n4434) );
  AND2X1 U4757 ( .A(\RF[0][41] ), .B(n10702), .Y(n2171) );
  INVX1 U4758 ( .A(n2171), .Y(n4435) );
  AND2X1 U4759 ( .A(\RF[0][29] ), .B(n10702), .Y(n2159) );
  INVX1 U4760 ( .A(n2159), .Y(n4436) );
  AND2X1 U4761 ( .A(\RF[0][17] ), .B(n10702), .Y(n2147) );
  INVX1 U4762 ( .A(n2147), .Y(n4437) );
  AND2X1 U4763 ( .A(\RF[0][5] ), .B(n10702), .Y(n2135) );
  INVX1 U4764 ( .A(n2135), .Y(n4438) );
  AND2X1 U4765 ( .A(\RF[1][38] ), .B(n10704), .Y(n2103) );
  INVX1 U4766 ( .A(n2103), .Y(n4439) );
  AND2X1 U4767 ( .A(\RF[1][30] ), .B(n10704), .Y(n2095) );
  INVX1 U4768 ( .A(n2095), .Y(n4440) );
  AND2X1 U4769 ( .A(\RF[1][18] ), .B(n10704), .Y(n2083) );
  INVX1 U4770 ( .A(n2083), .Y(n4441) );
  AND2X1 U4771 ( .A(\RF[1][6] ), .B(n10704), .Y(n2071) );
  INVX1 U4772 ( .A(n2071), .Y(n4442) );
  AND2X1 U4773 ( .A(\RF[2][43] ), .B(n10706), .Y(n2043) );
  INVX1 U4774 ( .A(n2043), .Y(n4443) );
  AND2X1 U4775 ( .A(\RF[2][31] ), .B(n10706), .Y(n2031) );
  INVX1 U4776 ( .A(n2031), .Y(n4444) );
  AND2X1 U4777 ( .A(\RF[2][19] ), .B(n10705), .Y(n2019) );
  INVX1 U4778 ( .A(n2019), .Y(n4445) );
  AND2X1 U4779 ( .A(\RF[2][7] ), .B(n10706), .Y(n2007) );
  INVX1 U4780 ( .A(n2007), .Y(n4446) );
  AND2X1 U4781 ( .A(\RF[3][47] ), .B(n10708), .Y(n1982) );
  INVX1 U4782 ( .A(n1982), .Y(n4447) );
  AND2X1 U4783 ( .A(\RF[3][25] ), .B(n10708), .Y(n1960) );
  INVX1 U4784 ( .A(n1960), .Y(n4448) );
  AND2X1 U4785 ( .A(\RF[3][20] ), .B(n10708), .Y(n1955) );
  INVX1 U4786 ( .A(n1955), .Y(n4449) );
  AND2X1 U4787 ( .A(\RF[3][8] ), .B(n10708), .Y(n1943) );
  INVX1 U4788 ( .A(n1943), .Y(n4450) );
  AND2X1 U4789 ( .A(\RF[4][44] ), .B(n10710), .Y(n1914) );
  INVX1 U4790 ( .A(n1914), .Y(n4451) );
  AND2X1 U4791 ( .A(\RF[4][33] ), .B(n10710), .Y(n1903) );
  INVX1 U4792 ( .A(n1903), .Y(n4452) );
  AND2X1 U4793 ( .A(\RF[4][21] ), .B(n10710), .Y(n1891) );
  INVX1 U4794 ( .A(n1891), .Y(n4453) );
  AND2X1 U4795 ( .A(\RF[4][9] ), .B(n10710), .Y(n1879) );
  INVX1 U4796 ( .A(n1879), .Y(n4454) );
  AND2X1 U4797 ( .A(\RF[5][63] ), .B(n10712), .Y(n1868) );
  INVX1 U4798 ( .A(n1868), .Y(n4455) );
  AND2X1 U4799 ( .A(\RF[5][34] ), .B(n10712), .Y(n1839) );
  INVX1 U4800 ( .A(n1839), .Y(n4456) );
  AND2X1 U4801 ( .A(\RF[5][22] ), .B(n10711), .Y(n1827) );
  INVX1 U4802 ( .A(n1827), .Y(n4457) );
  AND2X1 U4803 ( .A(\RF[5][10] ), .B(n10712), .Y(n1815) );
  INVX1 U4804 ( .A(n1815), .Y(n4458) );
  AND2X1 U4805 ( .A(\RF[6][56] ), .B(n10714), .Y(n1796) );
  INVX1 U4806 ( .A(n1796), .Y(n4459) );
  AND2X1 U4807 ( .A(\RF[6][35] ), .B(n10714), .Y(n1775) );
  INVX1 U4808 ( .A(n1775), .Y(n4460) );
  AND2X1 U4809 ( .A(\RF[6][23] ), .B(n10714), .Y(n1763) );
  INVX1 U4810 ( .A(n1763), .Y(n4461) );
  AND2X1 U4811 ( .A(\RF[6][11] ), .B(n10713), .Y(n1751) );
  INVX1 U4812 ( .A(n1751), .Y(n4462) );
  AND2X1 U4813 ( .A(\RF[7][59] ), .B(n10716), .Y(n1733) );
  INVX1 U4814 ( .A(n1733), .Y(n4463) );
  AND2X1 U4815 ( .A(\RF[7][42] ), .B(n10716), .Y(n1716) );
  INVX1 U4816 ( .A(n1716), .Y(n4464) );
  AND2X1 U4817 ( .A(\RF[7][36] ), .B(n10716), .Y(n1710) );
  INVX1 U4818 ( .A(n1710), .Y(n4465) );
  AND2X1 U4819 ( .A(\RF[7][12] ), .B(n10715), .Y(n1686) );
  INVX1 U4820 ( .A(n1686), .Y(n4466) );
  AND2X1 U4821 ( .A(\RF[8][57] ), .B(n10718), .Y(n1666) );
  INVX1 U4822 ( .A(n1666), .Y(n4467) );
  AND2X1 U4823 ( .A(\RF[8][46] ), .B(n10718), .Y(n1655) );
  INVX1 U4824 ( .A(n1655), .Y(n4468) );
  AND2X1 U4825 ( .A(\RF[8][24] ), .B(n10717), .Y(n1633) );
  INVX1 U4826 ( .A(n1633), .Y(n4469) );
  AND2X1 U4827 ( .A(\RF[9][58] ), .B(n10720), .Y(n1602) );
  INVX1 U4828 ( .A(n1602), .Y(n4470) );
  AND2X1 U4829 ( .A(\RF[9][48] ), .B(n10720), .Y(n1592) );
  INVX1 U4830 ( .A(n1592), .Y(n4471) );
  AND2X1 U4831 ( .A(\RF[10][61] ), .B(n10722), .Y(n1540) );
  INVX1 U4832 ( .A(n1540), .Y(n4472) );
  AND2X1 U4833 ( .A(\RF[10][53] ), .B(n10722), .Y(n1532) );
  INVX1 U4834 ( .A(n1532), .Y(n4473) );
  AND2X1 U4835 ( .A(\RF[10][49] ), .B(n10721), .Y(n1528) );
  INVX1 U4836 ( .A(n1528), .Y(n4474) );
  AND2X1 U4837 ( .A(\RF[11][50] ), .B(n10724), .Y(n1464) );
  INVX1 U4838 ( .A(n1464), .Y(n4475) );
  AND2X1 U4839 ( .A(\RF[12][41] ), .B(n10726), .Y(n1390) );
  INVX1 U4840 ( .A(n1390), .Y(n4476) );
  AND2X1 U4841 ( .A(\RF[12][29] ), .B(n10726), .Y(n1378) );
  INVX1 U4842 ( .A(n1378), .Y(n4477) );
  AND2X1 U4843 ( .A(\RF[12][17] ), .B(n10726), .Y(n1366) );
  INVX1 U4844 ( .A(n1366), .Y(n4478) );
  AND2X1 U4845 ( .A(\RF[12][5] ), .B(n10726), .Y(n1354) );
  INVX1 U4846 ( .A(n1354), .Y(n4479) );
  AND2X1 U4847 ( .A(\RF[13][38] ), .B(n10728), .Y(n1322) );
  INVX1 U4848 ( .A(n1322), .Y(n4480) );
  AND2X1 U4849 ( .A(\RF[13][30] ), .B(n10728), .Y(n1314) );
  INVX1 U4850 ( .A(n1314), .Y(n4481) );
  AND2X1 U4851 ( .A(\RF[13][18] ), .B(n10728), .Y(n1302) );
  INVX1 U4852 ( .A(n1302), .Y(n4482) );
  AND2X1 U4853 ( .A(\RF[13][6] ), .B(n10728), .Y(n1290) );
  INVX1 U4854 ( .A(n1290), .Y(n4483) );
  AND2X1 U4855 ( .A(\RF[14][43] ), .B(n10730), .Y(n1262) );
  INVX1 U4856 ( .A(n1262), .Y(n4484) );
  AND2X1 U4857 ( .A(\RF[14][31] ), .B(n10730), .Y(n1250) );
  INVX1 U4858 ( .A(n1250), .Y(n4485) );
  AND2X1 U4859 ( .A(\RF[14][19] ), .B(n10729), .Y(n1238) );
  INVX1 U4860 ( .A(n1238), .Y(n4486) );
  AND2X1 U4861 ( .A(\RF[14][7] ), .B(n10730), .Y(n1226) );
  INVX1 U4862 ( .A(n1226), .Y(n4487) );
  AND2X1 U4863 ( .A(\RF[15][47] ), .B(n10732), .Y(n1200) );
  INVX1 U4864 ( .A(n1200), .Y(n4488) );
  AND2X1 U4865 ( .A(\RF[15][25] ), .B(n10732), .Y(n1178) );
  INVX1 U4866 ( .A(n1178), .Y(n4489) );
  AND2X1 U4867 ( .A(\RF[15][20] ), .B(n10732), .Y(n1173) );
  INVX1 U4868 ( .A(n1173), .Y(n4490) );
  AND2X1 U4869 ( .A(\RF[15][8] ), .B(n10732), .Y(n1161) );
  INVX1 U4870 ( .A(n1161), .Y(n4491) );
  AND2X1 U4871 ( .A(\RF[16][44] ), .B(n10734), .Y(n1132) );
  INVX1 U4872 ( .A(n1132), .Y(n4492) );
  AND2X1 U4873 ( .A(\RF[16][33] ), .B(n10734), .Y(n1121) );
  INVX1 U4874 ( .A(n1121), .Y(n4493) );
  AND2X1 U4875 ( .A(\RF[16][21] ), .B(n10734), .Y(n1109) );
  INVX1 U4876 ( .A(n1109), .Y(n4494) );
  AND2X1 U4877 ( .A(\RF[16][9] ), .B(n10734), .Y(n1097) );
  INVX1 U4878 ( .A(n1097), .Y(n4495) );
  AND2X1 U4879 ( .A(\RF[17][63] ), .B(n10736), .Y(n1086) );
  INVX1 U4880 ( .A(n1086), .Y(n4496) );
  AND2X1 U4881 ( .A(\RF[17][34] ), .B(n10736), .Y(n1057) );
  INVX1 U4882 ( .A(n1057), .Y(n4497) );
  AND2X1 U4883 ( .A(\RF[17][22] ), .B(n10735), .Y(n1045) );
  INVX1 U4884 ( .A(n1045), .Y(n4498) );
  AND2X1 U4885 ( .A(\RF[17][10] ), .B(n10736), .Y(n1033) );
  INVX1 U4886 ( .A(n1033), .Y(n4499) );
  AND2X1 U4887 ( .A(\RF[18][56] ), .B(n10738), .Y(n1014) );
  INVX1 U4888 ( .A(n1014), .Y(n4500) );
  AND2X1 U4889 ( .A(\RF[18][35] ), .B(n10738), .Y(n993) );
  INVX1 U4890 ( .A(n993), .Y(n4501) );
  AND2X1 U4891 ( .A(\RF[18][23] ), .B(n10738), .Y(n981) );
  INVX1 U4892 ( .A(n981), .Y(n4502) );
  AND2X1 U4893 ( .A(\RF[18][11] ), .B(n10737), .Y(n969) );
  INVX1 U4894 ( .A(n969), .Y(n4503) );
  AND2X1 U4895 ( .A(\RF[19][59] ), .B(n10740), .Y(n952) );
  INVX1 U4896 ( .A(n952), .Y(n4504) );
  AND2X1 U4897 ( .A(\RF[19][42] ), .B(n10740), .Y(n935) );
  INVX1 U4898 ( .A(n935), .Y(n4505) );
  AND2X1 U4899 ( .A(\RF[19][36] ), .B(n10740), .Y(n929) );
  INVX1 U4900 ( .A(n929), .Y(n4506) );
  AND2X1 U4901 ( .A(\RF[19][12] ), .B(n10739), .Y(n905) );
  INVX1 U4902 ( .A(n905), .Y(n4507) );
  AND2X1 U4903 ( .A(\RF[20][57] ), .B(n10742), .Y(n885) );
  INVX1 U4904 ( .A(n885), .Y(n4508) );
  AND2X1 U4905 ( .A(\RF[20][46] ), .B(n10742), .Y(n874) );
  INVX1 U4906 ( .A(n874), .Y(n4509) );
  AND2X1 U4907 ( .A(\RF[20][24] ), .B(n10741), .Y(n852) );
  INVX1 U4908 ( .A(n852), .Y(n4510) );
  AND2X1 U4909 ( .A(\RF[21][58] ), .B(n10744), .Y(n821) );
  INVX1 U4910 ( .A(n821), .Y(n4511) );
  AND2X1 U4911 ( .A(\RF[21][48] ), .B(n10744), .Y(n811) );
  INVX1 U4912 ( .A(n811), .Y(n4512) );
  AND2X1 U4913 ( .A(\RF[22][61] ), .B(n10746), .Y(n759) );
  INVX1 U4914 ( .A(n759), .Y(n4513) );
  AND2X1 U4915 ( .A(\RF[22][53] ), .B(n10746), .Y(n751) );
  INVX1 U4916 ( .A(n751), .Y(n4514) );
  AND2X1 U4917 ( .A(\RF[22][49] ), .B(n10745), .Y(n747) );
  INVX1 U4918 ( .A(n747), .Y(n4515) );
  AND2X1 U4919 ( .A(\RF[23][50] ), .B(n10748), .Y(n682) );
  INVX1 U4920 ( .A(n682), .Y(n4516) );
  AND2X1 U4921 ( .A(\RF[24][44] ), .B(n10750), .Y(n609) );
  INVX1 U4922 ( .A(n609), .Y(n4517) );
  AND2X1 U4923 ( .A(\RF[24][33] ), .B(n10750), .Y(n598) );
  INVX1 U4924 ( .A(n598), .Y(n4518) );
  AND2X1 U4925 ( .A(\RF[24][21] ), .B(n10750), .Y(n586) );
  INVX1 U4926 ( .A(n586), .Y(n4519) );
  AND2X1 U4927 ( .A(\RF[24][9] ), .B(n10750), .Y(n574) );
  INVX1 U4928 ( .A(n574), .Y(n4520) );
  AND2X1 U4929 ( .A(\RF[25][63] ), .B(n10752), .Y(n562) );
  INVX1 U4930 ( .A(n562), .Y(n4521) );
  AND2X1 U4931 ( .A(\RF[25][34] ), .B(n10752), .Y(n533) );
  INVX1 U4932 ( .A(n533), .Y(n4522) );
  AND2X1 U4933 ( .A(\RF[25][22] ), .B(n10751), .Y(n521) );
  INVX1 U4934 ( .A(n521), .Y(n4523) );
  AND2X1 U4935 ( .A(\RF[25][10] ), .B(n10752), .Y(n509) );
  INVX1 U4936 ( .A(n509), .Y(n4524) );
  AND2X1 U4937 ( .A(\RF[26][56] ), .B(n10754), .Y(n489) );
  INVX1 U4938 ( .A(n489), .Y(n4525) );
  AND2X1 U4939 ( .A(\RF[26][35] ), .B(n10754), .Y(n468) );
  INVX1 U4940 ( .A(n468), .Y(n4526) );
  AND2X1 U4941 ( .A(\RF[26][23] ), .B(n10754), .Y(n456) );
  INVX1 U4942 ( .A(n456), .Y(n4527) );
  AND2X1 U4943 ( .A(\RF[26][11] ), .B(n10753), .Y(n444) );
  INVX1 U4944 ( .A(n444), .Y(n4528) );
  AND2X1 U4945 ( .A(\RF[27][59] ), .B(n10756), .Y(n426) );
  INVX1 U4946 ( .A(n426), .Y(n4529) );
  AND2X1 U4947 ( .A(\RF[27][42] ), .B(n10756), .Y(n409) );
  INVX1 U4948 ( .A(n409), .Y(n4530) );
  AND2X1 U4949 ( .A(\RF[27][36] ), .B(n10756), .Y(n403) );
  INVX1 U4950 ( .A(n403), .Y(n4531) );
  AND2X1 U4951 ( .A(\RF[27][12] ), .B(n10755), .Y(n379) );
  INVX1 U4952 ( .A(n379), .Y(n4532) );
  AND2X1 U4953 ( .A(\RF[28][57] ), .B(n10758), .Y(n358) );
  INVX1 U4954 ( .A(n358), .Y(n4533) );
  AND2X1 U4955 ( .A(\RF[28][46] ), .B(n10758), .Y(n347) );
  INVX1 U4956 ( .A(n347), .Y(n4534) );
  AND2X1 U4957 ( .A(\RF[28][24] ), .B(n10757), .Y(n325) );
  INVX1 U4958 ( .A(n325), .Y(n4535) );
  AND2X1 U4959 ( .A(\RF[29][58] ), .B(n10760), .Y(n293) );
  INVX1 U4960 ( .A(n293), .Y(n4536) );
  AND2X1 U4961 ( .A(\RF[29][48] ), .B(n10760), .Y(n283) );
  INVX1 U4962 ( .A(n283), .Y(n4537) );
  AND2X1 U4963 ( .A(\RF[30][61] ), .B(n10762), .Y(n230) );
  INVX1 U4964 ( .A(n230), .Y(n4538) );
  AND2X1 U4965 ( .A(\RF[30][53] ), .B(n10762), .Y(n222) );
  INVX1 U4966 ( .A(n222), .Y(n4539) );
  AND2X1 U4967 ( .A(\RF[30][49] ), .B(n10761), .Y(n218) );
  INVX1 U4968 ( .A(n218), .Y(n4540) );
  AND2X1 U4969 ( .A(\RF[31][50] ), .B(n10764), .Y(n139) );
  INVX1 U4970 ( .A(n139), .Y(n4541) );
  AND2X1 U4971 ( .A(\RF[0][38] ), .B(n10702), .Y(n2168) );
  INVX1 U4972 ( .A(n2168), .Y(n4542) );
  AND2X1 U4973 ( .A(\RF[0][30] ), .B(n10701), .Y(n2160) );
  INVX1 U4974 ( .A(n2160), .Y(n4543) );
  AND2X1 U4975 ( .A(\RF[0][18] ), .B(n10701), .Y(n2148) );
  INVX1 U4976 ( .A(n2148), .Y(n4544) );
  AND2X1 U4977 ( .A(\RF[0][6] ), .B(n10702), .Y(n2136) );
  INVX1 U4978 ( .A(n2136), .Y(n4545) );
  AND2X1 U4979 ( .A(\RF[1][41] ), .B(n10703), .Y(n2106) );
  INVX1 U4980 ( .A(n2106), .Y(n4546) );
  AND2X1 U4981 ( .A(\RF[1][29] ), .B(n10704), .Y(n2094) );
  INVX1 U4982 ( .A(n2094), .Y(n4547) );
  AND2X1 U4983 ( .A(\RF[1][17] ), .B(n10703), .Y(n2082) );
  INVX1 U4984 ( .A(n2082), .Y(n4548) );
  AND2X1 U4985 ( .A(\RF[1][5] ), .B(n10704), .Y(n2070) );
  INVX1 U4986 ( .A(n2070), .Y(n4549) );
  AND2X1 U4987 ( .A(\RF[2][47] ), .B(n10705), .Y(n2047) );
  INVX1 U4988 ( .A(n2047), .Y(n4550) );
  AND2X1 U4989 ( .A(\RF[2][25] ), .B(n10706), .Y(n2025) );
  INVX1 U4990 ( .A(n2025), .Y(n4551) );
  AND2X1 U4991 ( .A(\RF[2][20] ), .B(n10706), .Y(n2020) );
  INVX1 U4992 ( .A(n2020), .Y(n4552) );
  AND2X1 U4993 ( .A(\RF[2][8] ), .B(n10706), .Y(n2008) );
  INVX1 U4994 ( .A(n2008), .Y(n4553) );
  AND2X1 U4995 ( .A(\RF[3][43] ), .B(n10707), .Y(n1978) );
  INVX1 U4996 ( .A(n1978), .Y(n4554) );
  AND2X1 U4997 ( .A(\RF[3][31] ), .B(n10708), .Y(n1966) );
  INVX1 U4998 ( .A(n1966), .Y(n4555) );
  AND2X1 U4999 ( .A(\RF[3][19] ), .B(n10708), .Y(n1954) );
  INVX1 U5000 ( .A(n1954), .Y(n4556) );
  AND2X1 U5001 ( .A(\RF[3][7] ), .B(n10708), .Y(n1942) );
  INVX1 U5002 ( .A(n1942), .Y(n4557) );
  AND2X1 U5003 ( .A(\RF[4][63] ), .B(n10710), .Y(n1933) );
  INVX1 U5004 ( .A(n1933), .Y(n4558) );
  AND2X1 U5005 ( .A(\RF[4][34] ), .B(n10710), .Y(n1904) );
  INVX1 U5006 ( .A(n1904), .Y(n4559) );
  AND2X1 U5007 ( .A(\RF[4][22] ), .B(n10710), .Y(n1892) );
  INVX1 U5008 ( .A(n1892), .Y(n4560) );
  AND2X1 U5009 ( .A(\RF[4][10] ), .B(n10710), .Y(n1880) );
  INVX1 U5010 ( .A(n1880), .Y(n4561) );
  AND2X1 U5011 ( .A(\RF[5][44] ), .B(n10712), .Y(n1849) );
  INVX1 U5012 ( .A(n1849), .Y(n4562) );
  AND2X1 U5013 ( .A(\RF[5][33] ), .B(n10712), .Y(n1838) );
  INVX1 U5014 ( .A(n1838), .Y(n4563) );
  AND2X1 U5015 ( .A(\RF[5][21] ), .B(n10712), .Y(n1826) );
  INVX1 U5016 ( .A(n1826), .Y(n4564) );
  AND2X1 U5017 ( .A(\RF[5][9] ), .B(n10712), .Y(n1814) );
  INVX1 U5018 ( .A(n1814), .Y(n4565) );
  AND2X1 U5019 ( .A(\RF[6][59] ), .B(n10714), .Y(n1799) );
  INVX1 U5020 ( .A(n1799), .Y(n4566) );
  AND2X1 U5021 ( .A(\RF[6][42] ), .B(n10714), .Y(n1782) );
  INVX1 U5022 ( .A(n1782), .Y(n4567) );
  AND2X1 U5023 ( .A(\RF[6][36] ), .B(n10713), .Y(n1776) );
  INVX1 U5024 ( .A(n1776), .Y(n4568) );
  AND2X1 U5025 ( .A(\RF[6][12] ), .B(n10714), .Y(n1752) );
  INVX1 U5026 ( .A(n1752), .Y(n4569) );
  AND2X1 U5027 ( .A(\RF[7][56] ), .B(n10716), .Y(n1730) );
  INVX1 U5028 ( .A(n1730), .Y(n4570) );
  AND2X1 U5029 ( .A(\RF[7][35] ), .B(n10715), .Y(n1709) );
  INVX1 U5030 ( .A(n1709), .Y(n4571) );
  AND2X1 U5031 ( .A(\RF[7][23] ), .B(n10716), .Y(n1697) );
  INVX1 U5032 ( .A(n1697), .Y(n4572) );
  AND2X1 U5033 ( .A(\RF[7][11] ), .B(n10716), .Y(n1685) );
  INVX1 U5034 ( .A(n1685), .Y(n4573) );
  AND2X1 U5035 ( .A(\RF[8][58] ), .B(n10718), .Y(n1667) );
  INVX1 U5036 ( .A(n1667), .Y(n4574) );
  AND2X1 U5037 ( .A(\RF[8][48] ), .B(n10718), .Y(n1657) );
  INVX1 U5038 ( .A(n1657), .Y(n4575) );
  AND2X1 U5039 ( .A(\RF[9][57] ), .B(n10720), .Y(n1601) );
  INVX1 U5040 ( .A(n1601), .Y(n4576) );
  AND2X1 U5041 ( .A(\RF[9][46] ), .B(n10720), .Y(n1590) );
  INVX1 U5042 ( .A(n1590), .Y(n4577) );
  AND2X1 U5043 ( .A(\RF[9][24] ), .B(n10719), .Y(n1568) );
  INVX1 U5044 ( .A(n1568), .Y(n4578) );
  AND2X1 U5045 ( .A(\RF[10][50] ), .B(n10722), .Y(n1529) );
  INVX1 U5046 ( .A(n1529), .Y(n4579) );
  AND2X1 U5047 ( .A(\RF[11][61] ), .B(n10724), .Y(n1475) );
  INVX1 U5048 ( .A(n1475), .Y(n4580) );
  AND2X1 U5049 ( .A(\RF[11][53] ), .B(n10724), .Y(n1467) );
  INVX1 U5050 ( .A(n1467), .Y(n4581) );
  AND2X1 U5051 ( .A(\RF[11][49] ), .B(n10723), .Y(n1463) );
  INVX1 U5052 ( .A(n1463), .Y(n4582) );
  AND2X1 U5053 ( .A(\RF[12][38] ), .B(n10726), .Y(n1387) );
  INVX1 U5054 ( .A(n1387), .Y(n4583) );
  AND2X1 U5055 ( .A(\RF[12][30] ), .B(n10725), .Y(n1379) );
  INVX1 U5056 ( .A(n1379), .Y(n4584) );
  AND2X1 U5057 ( .A(\RF[12][18] ), .B(n10725), .Y(n1367) );
  INVX1 U5058 ( .A(n1367), .Y(n4585) );
  AND2X1 U5059 ( .A(\RF[12][6] ), .B(n10726), .Y(n1355) );
  INVX1 U5060 ( .A(n1355), .Y(n4586) );
  AND2X1 U5061 ( .A(\RF[13][41] ), .B(n10727), .Y(n1325) );
  INVX1 U5062 ( .A(n1325), .Y(n4587) );
  AND2X1 U5063 ( .A(\RF[13][29] ), .B(n10728), .Y(n1313) );
  INVX1 U5064 ( .A(n1313), .Y(n4588) );
  AND2X1 U5065 ( .A(\RF[13][17] ), .B(n10727), .Y(n1301) );
  INVX1 U5066 ( .A(n1301), .Y(n4589) );
  AND2X1 U5067 ( .A(\RF[13][5] ), .B(n10728), .Y(n1289) );
  INVX1 U5068 ( .A(n1289), .Y(n4590) );
  AND2X1 U5069 ( .A(\RF[14][47] ), .B(n10729), .Y(n1266) );
  INVX1 U5070 ( .A(n1266), .Y(n4591) );
  AND2X1 U5071 ( .A(\RF[14][25] ), .B(n10730), .Y(n1244) );
  INVX1 U5072 ( .A(n1244), .Y(n4592) );
  AND2X1 U5073 ( .A(\RF[14][20] ), .B(n10730), .Y(n1239) );
  INVX1 U5074 ( .A(n1239), .Y(n4593) );
  AND2X1 U5075 ( .A(\RF[14][8] ), .B(n10730), .Y(n1227) );
  INVX1 U5076 ( .A(n1227), .Y(n4594) );
  AND2X1 U5077 ( .A(\RF[15][43] ), .B(n10731), .Y(n1196) );
  INVX1 U5078 ( .A(n1196), .Y(n4595) );
  AND2X1 U5079 ( .A(\RF[15][31] ), .B(n10732), .Y(n1184) );
  INVX1 U5080 ( .A(n1184), .Y(n4596) );
  AND2X1 U5081 ( .A(\RF[15][19] ), .B(n10732), .Y(n1172) );
  INVX1 U5082 ( .A(n1172), .Y(n4597) );
  AND2X1 U5083 ( .A(\RF[15][7] ), .B(n10732), .Y(n1160) );
  INVX1 U5084 ( .A(n1160), .Y(n4598) );
  AND2X1 U5085 ( .A(\RF[16][63] ), .B(n10734), .Y(n1151) );
  INVX1 U5086 ( .A(n1151), .Y(n4599) );
  AND2X1 U5087 ( .A(\RF[16][34] ), .B(n10734), .Y(n1122) );
  INVX1 U5088 ( .A(n1122), .Y(n4600) );
  AND2X1 U5089 ( .A(\RF[16][22] ), .B(n10734), .Y(n1110) );
  INVX1 U5090 ( .A(n1110), .Y(n4601) );
  AND2X1 U5091 ( .A(\RF[16][10] ), .B(n10734), .Y(n1098) );
  INVX1 U5092 ( .A(n1098), .Y(n4602) );
  AND2X1 U5093 ( .A(\RF[17][44] ), .B(n10736), .Y(n1067) );
  INVX1 U5094 ( .A(n1067), .Y(n4603) );
  AND2X1 U5095 ( .A(\RF[17][33] ), .B(n10736), .Y(n1056) );
  INVX1 U5096 ( .A(n1056), .Y(n4604) );
  AND2X1 U5097 ( .A(\RF[17][21] ), .B(n10736), .Y(n1044) );
  INVX1 U5098 ( .A(n1044), .Y(n4605) );
  AND2X1 U5099 ( .A(\RF[17][9] ), .B(n10736), .Y(n1032) );
  INVX1 U5100 ( .A(n1032), .Y(n4606) );
  AND2X1 U5101 ( .A(\RF[18][59] ), .B(n10738), .Y(n1017) );
  INVX1 U5102 ( .A(n1017), .Y(n4607) );
  AND2X1 U5103 ( .A(\RF[18][42] ), .B(n10738), .Y(n1000) );
  INVX1 U5104 ( .A(n1000), .Y(n4608) );
  AND2X1 U5105 ( .A(\RF[18][36] ), .B(n10737), .Y(n994) );
  INVX1 U5106 ( .A(n994), .Y(n4609) );
  AND2X1 U5107 ( .A(\RF[18][12] ), .B(n10738), .Y(n970) );
  INVX1 U5108 ( .A(n970), .Y(n4610) );
  AND2X1 U5109 ( .A(\RF[19][56] ), .B(n10740), .Y(n949) );
  INVX1 U5110 ( .A(n949), .Y(n4611) );
  AND2X1 U5111 ( .A(\RF[19][35] ), .B(n10739), .Y(n928) );
  INVX1 U5112 ( .A(n928), .Y(n4612) );
  AND2X1 U5113 ( .A(\RF[19][23] ), .B(n10740), .Y(n916) );
  INVX1 U5114 ( .A(n916), .Y(n4613) );
  AND2X1 U5115 ( .A(\RF[19][11] ), .B(n10740), .Y(n904) );
  INVX1 U5116 ( .A(n904), .Y(n4614) );
  AND2X1 U5117 ( .A(\RF[20][58] ), .B(n10742), .Y(n886) );
  INVX1 U5118 ( .A(n886), .Y(n4615) );
  AND2X1 U5119 ( .A(\RF[20][48] ), .B(n10742), .Y(n876) );
  INVX1 U5120 ( .A(n876), .Y(n4616) );
  AND2X1 U5121 ( .A(\RF[21][57] ), .B(n10744), .Y(n820) );
  INVX1 U5122 ( .A(n820), .Y(n4617) );
  AND2X1 U5123 ( .A(\RF[21][46] ), .B(n10744), .Y(n809) );
  INVX1 U5124 ( .A(n809), .Y(n4618) );
  AND2X1 U5125 ( .A(\RF[21][24] ), .B(n10743), .Y(n787) );
  INVX1 U5126 ( .A(n787), .Y(n4619) );
  AND2X1 U5127 ( .A(\RF[22][50] ), .B(n10746), .Y(n748) );
  INVX1 U5128 ( .A(n748), .Y(n4620) );
  AND2X1 U5129 ( .A(\RF[23][61] ), .B(n10748), .Y(n693) );
  INVX1 U5130 ( .A(n693), .Y(n4621) );
  AND2X1 U5131 ( .A(\RF[23][53] ), .B(n10748), .Y(n685) );
  INVX1 U5132 ( .A(n685), .Y(n4622) );
  AND2X1 U5133 ( .A(\RF[23][49] ), .B(n10747), .Y(n681) );
  INVX1 U5134 ( .A(n681), .Y(n4623) );
  AND2X1 U5135 ( .A(\RF[24][63] ), .B(n10750), .Y(n628) );
  INVX1 U5136 ( .A(n628), .Y(n4624) );
  AND2X1 U5137 ( .A(\RF[24][34] ), .B(n10750), .Y(n599) );
  INVX1 U5138 ( .A(n599), .Y(n4625) );
  AND2X1 U5139 ( .A(\RF[24][22] ), .B(n10750), .Y(n587) );
  INVX1 U5140 ( .A(n587), .Y(n4626) );
  AND2X1 U5141 ( .A(\RF[24][10] ), .B(n10750), .Y(n575) );
  INVX1 U5142 ( .A(n575), .Y(n4627) );
  AND2X1 U5143 ( .A(\RF[25][44] ), .B(n10752), .Y(n543) );
  INVX1 U5144 ( .A(n543), .Y(n4628) );
  AND2X1 U5145 ( .A(\RF[25][33] ), .B(n10752), .Y(n532) );
  INVX1 U5146 ( .A(n532), .Y(n4629) );
  AND2X1 U5147 ( .A(\RF[25][21] ), .B(n10752), .Y(n520) );
  INVX1 U5148 ( .A(n520), .Y(n4630) );
  AND2X1 U5149 ( .A(\RF[25][9] ), .B(n10752), .Y(n508) );
  INVX1 U5150 ( .A(n508), .Y(n4631) );
  AND2X1 U5151 ( .A(\RF[26][59] ), .B(n10754), .Y(n492) );
  INVX1 U5152 ( .A(n492), .Y(n4632) );
  AND2X1 U5153 ( .A(\RF[26][42] ), .B(n10754), .Y(n475) );
  INVX1 U5154 ( .A(n475), .Y(n4633) );
  AND2X1 U5155 ( .A(\RF[26][36] ), .B(n10753), .Y(n469) );
  INVX1 U5156 ( .A(n469), .Y(n4634) );
  AND2X1 U5157 ( .A(\RF[26][12] ), .B(n10754), .Y(n445) );
  INVX1 U5158 ( .A(n445), .Y(n4635) );
  AND2X1 U5159 ( .A(\RF[27][56] ), .B(n10756), .Y(n423) );
  INVX1 U5160 ( .A(n423), .Y(n4636) );
  AND2X1 U5161 ( .A(\RF[27][35] ), .B(n10755), .Y(n402) );
  INVX1 U5162 ( .A(n402), .Y(n4637) );
  AND2X1 U5163 ( .A(\RF[27][23] ), .B(n10756), .Y(n390) );
  INVX1 U5164 ( .A(n390), .Y(n4638) );
  AND2X1 U5165 ( .A(\RF[27][11] ), .B(n10756), .Y(n378) );
  INVX1 U5166 ( .A(n378), .Y(n4639) );
  AND2X1 U5167 ( .A(\RF[28][58] ), .B(n10758), .Y(n359) );
  INVX1 U5168 ( .A(n359), .Y(n4640) );
  AND2X1 U5169 ( .A(\RF[28][48] ), .B(n10758), .Y(n349) );
  INVX1 U5170 ( .A(n349), .Y(n4641) );
  AND2X1 U5171 ( .A(\RF[29][57] ), .B(n10760), .Y(n292) );
  INVX1 U5172 ( .A(n292), .Y(n4642) );
  AND2X1 U5173 ( .A(\RF[29][46] ), .B(n10760), .Y(n281) );
  INVX1 U5174 ( .A(n281), .Y(n4643) );
  AND2X1 U5175 ( .A(\RF[29][24] ), .B(n10759), .Y(n259) );
  INVX1 U5176 ( .A(n259), .Y(n4644) );
  AND2X1 U5177 ( .A(\RF[30][50] ), .B(n10762), .Y(n219) );
  INVX1 U5178 ( .A(n219), .Y(n4645) );
  AND2X1 U5179 ( .A(\RF[31][61] ), .B(n10764), .Y(n161) );
  INVX1 U5180 ( .A(n161), .Y(n4646) );
  AND2X1 U5181 ( .A(\RF[31][53] ), .B(n10764), .Y(n145) );
  INVX1 U5182 ( .A(n145), .Y(n4647) );
  AND2X1 U5183 ( .A(\RF[31][49] ), .B(n10763), .Y(n137) );
  INVX1 U5184 ( .A(n137), .Y(n4648) );
  AND2X1 U5185 ( .A(\RF[0][43] ), .B(n10702), .Y(n2173) );
  INVX1 U5186 ( .A(n2173), .Y(n4649) );
  AND2X1 U5187 ( .A(\RF[0][31] ), .B(n10701), .Y(n2161) );
  INVX1 U5188 ( .A(n2161), .Y(n4650) );
  AND2X1 U5189 ( .A(\RF[0][19] ), .B(n10702), .Y(n2149) );
  INVX1 U5190 ( .A(n2149), .Y(n4651) );
  AND2X1 U5191 ( .A(\RF[0][7] ), .B(n10702), .Y(n2137) );
  INVX1 U5192 ( .A(n2137), .Y(n4652) );
  AND2X1 U5193 ( .A(\RF[1][47] ), .B(n10704), .Y(n2112) );
  INVX1 U5194 ( .A(n2112), .Y(n4653) );
  AND2X1 U5195 ( .A(\RF[1][25] ), .B(n10704), .Y(n2090) );
  INVX1 U5196 ( .A(n2090), .Y(n4654) );
  AND2X1 U5197 ( .A(\RF[1][20] ), .B(n10703), .Y(n2085) );
  INVX1 U5198 ( .A(n2085), .Y(n4655) );
  AND2X1 U5199 ( .A(\RF[1][8] ), .B(n10704), .Y(n2073) );
  INVX1 U5200 ( .A(n2073), .Y(n4656) );
  AND2X1 U5201 ( .A(\RF[2][41] ), .B(n10706), .Y(n2041) );
  INVX1 U5202 ( .A(n2041), .Y(n4657) );
  AND2X1 U5203 ( .A(\RF[2][29] ), .B(n10706), .Y(n2029) );
  INVX1 U5204 ( .A(n2029), .Y(n4658) );
  AND2X1 U5205 ( .A(\RF[2][17] ), .B(n10705), .Y(n2017) );
  INVX1 U5206 ( .A(n2017), .Y(n4659) );
  AND2X1 U5207 ( .A(\RF[2][5] ), .B(n10705), .Y(n2005) );
  INVX1 U5208 ( .A(n2005), .Y(n4660) );
  AND2X1 U5209 ( .A(\RF[3][38] ), .B(n10707), .Y(n1973) );
  INVX1 U5210 ( .A(n1973), .Y(n4661) );
  AND2X1 U5211 ( .A(\RF[3][30] ), .B(n10708), .Y(n1965) );
  INVX1 U5212 ( .A(n1965), .Y(n4662) );
  AND2X1 U5213 ( .A(\RF[3][18] ), .B(n10708), .Y(n1953) );
  INVX1 U5214 ( .A(n1953), .Y(n4663) );
  AND2X1 U5215 ( .A(\RF[3][6] ), .B(n10707), .Y(n1941) );
  INVX1 U5216 ( .A(n1941), .Y(n4664) );
  AND2X1 U5217 ( .A(\RF[4][56] ), .B(n10709), .Y(n1926) );
  INVX1 U5218 ( .A(n1926), .Y(n4665) );
  AND2X1 U5219 ( .A(\RF[4][35] ), .B(n10709), .Y(n1905) );
  INVX1 U5220 ( .A(n1905), .Y(n4666) );
  AND2X1 U5221 ( .A(\RF[4][23] ), .B(n10709), .Y(n1893) );
  INVX1 U5222 ( .A(n1893), .Y(n4667) );
  AND2X1 U5223 ( .A(\RF[4][11] ), .B(n10710), .Y(n1881) );
  INVX1 U5224 ( .A(n1881), .Y(n4668) );
  AND2X1 U5225 ( .A(\RF[5][59] ), .B(n10711), .Y(n1864) );
  INVX1 U5226 ( .A(n1864), .Y(n4669) );
  AND2X1 U5227 ( .A(\RF[5][42] ), .B(n10712), .Y(n1847) );
  INVX1 U5228 ( .A(n1847), .Y(n4670) );
  AND2X1 U5229 ( .A(\RF[5][36] ), .B(n10711), .Y(n1841) );
  INVX1 U5230 ( .A(n1841), .Y(n4671) );
  AND2X1 U5231 ( .A(\RF[5][12] ), .B(n10711), .Y(n1817) );
  INVX1 U5232 ( .A(n1817), .Y(n4672) );
  AND2X1 U5233 ( .A(\RF[6][44] ), .B(n10713), .Y(n1784) );
  INVX1 U5234 ( .A(n1784), .Y(n4673) );
  AND2X1 U5235 ( .A(\RF[6][33] ), .B(n10714), .Y(n1773) );
  INVX1 U5236 ( .A(n1773), .Y(n4674) );
  AND2X1 U5237 ( .A(\RF[6][21] ), .B(n10714), .Y(n1761) );
  INVX1 U5238 ( .A(n1761), .Y(n4675) );
  AND2X1 U5239 ( .A(\RF[6][9] ), .B(n10713), .Y(n1749) );
  INVX1 U5240 ( .A(n1749), .Y(n4676) );
  AND2X1 U5241 ( .A(\RF[7][63] ), .B(n10716), .Y(n1737) );
  INVX1 U5242 ( .A(n1737), .Y(n4677) );
  AND2X1 U5243 ( .A(\RF[7][34] ), .B(n10716), .Y(n1708) );
  INVX1 U5244 ( .A(n1708), .Y(n4678) );
  AND2X1 U5245 ( .A(\RF[7][22] ), .B(n10715), .Y(n1696) );
  INVX1 U5246 ( .A(n1696), .Y(n4679) );
  AND2X1 U5247 ( .A(\RF[7][10] ), .B(n10715), .Y(n1684) );
  INVX1 U5248 ( .A(n1684), .Y(n4680) );
  AND2X1 U5249 ( .A(\RF[8][61] ), .B(n10717), .Y(n1670) );
  INVX1 U5250 ( .A(n1670), .Y(n4681) );
  AND2X1 U5251 ( .A(\RF[8][53] ), .B(n10718), .Y(n1662) );
  INVX1 U5252 ( .A(n1662), .Y(n4682) );
  AND2X1 U5253 ( .A(\RF[8][49] ), .B(n10718), .Y(n1658) );
  INVX1 U5254 ( .A(n1658), .Y(n4683) );
  AND2X1 U5255 ( .A(\RF[9][50] ), .B(n10720), .Y(n1594) );
  INVX1 U5256 ( .A(n1594), .Y(n4684) );
  AND2X1 U5257 ( .A(\RF[10][57] ), .B(n10722), .Y(n1536) );
  INVX1 U5258 ( .A(n1536), .Y(n4685) );
  AND2X1 U5259 ( .A(\RF[10][46] ), .B(n10722), .Y(n1525) );
  INVX1 U5260 ( .A(n1525), .Y(n4686) );
  AND2X1 U5261 ( .A(\RF[10][24] ), .B(n10722), .Y(n1503) );
  INVX1 U5262 ( .A(n1503), .Y(n4687) );
  AND2X1 U5263 ( .A(\RF[11][58] ), .B(n10724), .Y(n1472) );
  INVX1 U5264 ( .A(n1472), .Y(n4688) );
  AND2X1 U5265 ( .A(\RF[11][48] ), .B(n10724), .Y(n1462) );
  INVX1 U5266 ( .A(n1462), .Y(n4689) );
  AND2X1 U5267 ( .A(\RF[12][43] ), .B(n10726), .Y(n1392) );
  INVX1 U5268 ( .A(n1392), .Y(n4690) );
  AND2X1 U5269 ( .A(\RF[12][31] ), .B(n10725), .Y(n1380) );
  INVX1 U5270 ( .A(n1380), .Y(n4691) );
  AND2X1 U5271 ( .A(\RF[12][19] ), .B(n10726), .Y(n1368) );
  INVX1 U5272 ( .A(n1368), .Y(n4692) );
  AND2X1 U5273 ( .A(\RF[12][7] ), .B(n10726), .Y(n1356) );
  INVX1 U5274 ( .A(n1356), .Y(n4693) );
  AND2X1 U5275 ( .A(\RF[13][47] ), .B(n10728), .Y(n1331) );
  INVX1 U5276 ( .A(n1331), .Y(n4694) );
  AND2X1 U5277 ( .A(\RF[13][25] ), .B(n10728), .Y(n1309) );
  INVX1 U5278 ( .A(n1309), .Y(n4695) );
  AND2X1 U5279 ( .A(\RF[13][20] ), .B(n10727), .Y(n1304) );
  INVX1 U5280 ( .A(n1304), .Y(n4696) );
  AND2X1 U5281 ( .A(\RF[13][8] ), .B(n10728), .Y(n1292) );
  INVX1 U5282 ( .A(n1292), .Y(n4697) );
  AND2X1 U5283 ( .A(\RF[14][41] ), .B(n10730), .Y(n1260) );
  INVX1 U5284 ( .A(n1260), .Y(n4698) );
  AND2X1 U5285 ( .A(\RF[14][29] ), .B(n10730), .Y(n1248) );
  INVX1 U5286 ( .A(n1248), .Y(n4699) );
  AND2X1 U5287 ( .A(\RF[14][17] ), .B(n10729), .Y(n1236) );
  INVX1 U5288 ( .A(n1236), .Y(n4700) );
  AND2X1 U5289 ( .A(\RF[14][5] ), .B(n10729), .Y(n1224) );
  INVX1 U5290 ( .A(n1224), .Y(n4701) );
  AND2X1 U5291 ( .A(\RF[15][38] ), .B(n10731), .Y(n1191) );
  INVX1 U5292 ( .A(n1191), .Y(n4702) );
  AND2X1 U5293 ( .A(\RF[15][30] ), .B(n10732), .Y(n1183) );
  INVX1 U5294 ( .A(n1183), .Y(n4703) );
  AND2X1 U5295 ( .A(\RF[15][18] ), .B(n10732), .Y(n1171) );
  INVX1 U5296 ( .A(n1171), .Y(n4704) );
  AND2X1 U5297 ( .A(\RF[15][6] ), .B(n10731), .Y(n1159) );
  INVX1 U5298 ( .A(n1159), .Y(n4705) );
  AND2X1 U5299 ( .A(\RF[16][56] ), .B(n10733), .Y(n1144) );
  INVX1 U5300 ( .A(n1144), .Y(n4706) );
  AND2X1 U5301 ( .A(\RF[16][35] ), .B(n10733), .Y(n1123) );
  INVX1 U5302 ( .A(n1123), .Y(n4707) );
  AND2X1 U5303 ( .A(\RF[16][23] ), .B(n10733), .Y(n1111) );
  INVX1 U5304 ( .A(n1111), .Y(n4708) );
  AND2X1 U5305 ( .A(\RF[16][11] ), .B(n10734), .Y(n1099) );
  INVX1 U5306 ( .A(n1099), .Y(n4709) );
  AND2X1 U5307 ( .A(\RF[17][59] ), .B(n10735), .Y(n1082) );
  INVX1 U5308 ( .A(n1082), .Y(n4710) );
  AND2X1 U5309 ( .A(\RF[17][42] ), .B(n10736), .Y(n1065) );
  INVX1 U5310 ( .A(n1065), .Y(n4711) );
  AND2X1 U5311 ( .A(\RF[17][36] ), .B(n10735), .Y(n1059) );
  INVX1 U5312 ( .A(n1059), .Y(n4712) );
  AND2X1 U5313 ( .A(\RF[17][12] ), .B(n10735), .Y(n1035) );
  INVX1 U5314 ( .A(n1035), .Y(n4713) );
  AND2X1 U5315 ( .A(\RF[18][44] ), .B(n10737), .Y(n1002) );
  INVX1 U5316 ( .A(n1002), .Y(n4714) );
  AND2X1 U5317 ( .A(\RF[18][33] ), .B(n10738), .Y(n991) );
  INVX1 U5318 ( .A(n991), .Y(n4715) );
  AND2X1 U5319 ( .A(\RF[18][21] ), .B(n10738), .Y(n979) );
  INVX1 U5320 ( .A(n979), .Y(n4716) );
  AND2X1 U5321 ( .A(\RF[18][9] ), .B(n10737), .Y(n967) );
  INVX1 U5322 ( .A(n967), .Y(n4717) );
  AND2X1 U5323 ( .A(\RF[19][63] ), .B(n10740), .Y(n956) );
  INVX1 U5324 ( .A(n956), .Y(n4718) );
  AND2X1 U5325 ( .A(\RF[19][34] ), .B(n10740), .Y(n927) );
  INVX1 U5326 ( .A(n927), .Y(n4719) );
  AND2X1 U5327 ( .A(\RF[19][22] ), .B(n10739), .Y(n915) );
  INVX1 U5328 ( .A(n915), .Y(n4720) );
  AND2X1 U5329 ( .A(\RF[19][10] ), .B(n10739), .Y(n903) );
  INVX1 U5330 ( .A(n903), .Y(n4721) );
  AND2X1 U5331 ( .A(\RF[20][61] ), .B(n10741), .Y(n889) );
  INVX1 U5332 ( .A(n889), .Y(n4722) );
  AND2X1 U5333 ( .A(\RF[20][53] ), .B(n10742), .Y(n881) );
  INVX1 U5334 ( .A(n881), .Y(n4723) );
  AND2X1 U5335 ( .A(\RF[20][49] ), .B(n10742), .Y(n877) );
  INVX1 U5336 ( .A(n877), .Y(n4724) );
  AND2X1 U5337 ( .A(\RF[21][50] ), .B(n10744), .Y(n813) );
  INVX1 U5338 ( .A(n813), .Y(n4725) );
  AND2X1 U5339 ( .A(\RF[22][57] ), .B(n10746), .Y(n755) );
  INVX1 U5340 ( .A(n755), .Y(n4726) );
  AND2X1 U5341 ( .A(\RF[22][46] ), .B(n10746), .Y(n744) );
  INVX1 U5342 ( .A(n744), .Y(n4727) );
  AND2X1 U5343 ( .A(\RF[22][24] ), .B(n10746), .Y(n722) );
  INVX1 U5344 ( .A(n722), .Y(n4728) );
  AND2X1 U5345 ( .A(\RF[23][58] ), .B(n10748), .Y(n690) );
  INVX1 U5346 ( .A(n690), .Y(n4729) );
  AND2X1 U5347 ( .A(\RF[23][48] ), .B(n10748), .Y(n680) );
  INVX1 U5348 ( .A(n680), .Y(n4730) );
  AND2X1 U5349 ( .A(\RF[24][56] ), .B(n10749), .Y(n621) );
  INVX1 U5350 ( .A(n621), .Y(n4731) );
  AND2X1 U5351 ( .A(\RF[24][35] ), .B(n10749), .Y(n600) );
  INVX1 U5352 ( .A(n600), .Y(n4732) );
  AND2X1 U5353 ( .A(\RF[24][23] ), .B(n10749), .Y(n588) );
  INVX1 U5354 ( .A(n588), .Y(n4733) );
  AND2X1 U5355 ( .A(\RF[24][11] ), .B(n10750), .Y(n576) );
  INVX1 U5356 ( .A(n576), .Y(n4734) );
  AND2X1 U5357 ( .A(\RF[25][59] ), .B(n10751), .Y(n558) );
  INVX1 U5358 ( .A(n558), .Y(n4735) );
  AND2X1 U5359 ( .A(\RF[25][42] ), .B(n10752), .Y(n541) );
  INVX1 U5360 ( .A(n541), .Y(n4736) );
  AND2X1 U5361 ( .A(\RF[25][36] ), .B(n10751), .Y(n535) );
  INVX1 U5362 ( .A(n535), .Y(n4737) );
  AND2X1 U5363 ( .A(\RF[25][12] ), .B(n10751), .Y(n511) );
  INVX1 U5364 ( .A(n511), .Y(n4738) );
  AND2X1 U5365 ( .A(\RF[26][44] ), .B(n10753), .Y(n477) );
  INVX1 U5366 ( .A(n477), .Y(n4739) );
  AND2X1 U5367 ( .A(\RF[26][33] ), .B(n10754), .Y(n466) );
  INVX1 U5368 ( .A(n466), .Y(n4740) );
  AND2X1 U5369 ( .A(\RF[26][21] ), .B(n10754), .Y(n454) );
  INVX1 U5370 ( .A(n454), .Y(n4741) );
  AND2X1 U5371 ( .A(\RF[26][9] ), .B(n10753), .Y(n442) );
  INVX1 U5372 ( .A(n442), .Y(n4742) );
  AND2X1 U5373 ( .A(\RF[27][63] ), .B(n10756), .Y(n430) );
  INVX1 U5374 ( .A(n430), .Y(n4743) );
  AND2X1 U5375 ( .A(\RF[27][34] ), .B(n10756), .Y(n401) );
  INVX1 U5376 ( .A(n401), .Y(n4744) );
  AND2X1 U5377 ( .A(\RF[27][22] ), .B(n10755), .Y(n389) );
  INVX1 U5378 ( .A(n389), .Y(n4745) );
  AND2X1 U5379 ( .A(\RF[27][10] ), .B(n10755), .Y(n377) );
  INVX1 U5380 ( .A(n377), .Y(n4746) );
  AND2X1 U5381 ( .A(\RF[28][61] ), .B(n10757), .Y(n362) );
  INVX1 U5382 ( .A(n362), .Y(n4747) );
  AND2X1 U5383 ( .A(\RF[28][53] ), .B(n10758), .Y(n354) );
  INVX1 U5384 ( .A(n354), .Y(n4748) );
  AND2X1 U5385 ( .A(\RF[28][49] ), .B(n10758), .Y(n350) );
  INVX1 U5386 ( .A(n350), .Y(n4749) );
  AND2X1 U5387 ( .A(\RF[29][50] ), .B(n10760), .Y(n285) );
  INVX1 U5388 ( .A(n285), .Y(n4750) );
  AND2X1 U5389 ( .A(\RF[30][57] ), .B(n10762), .Y(n226) );
  INVX1 U5390 ( .A(n226), .Y(n4751) );
  AND2X1 U5391 ( .A(\RF[30][46] ), .B(n10762), .Y(n215) );
  INVX1 U5392 ( .A(n215), .Y(n4752) );
  AND2X1 U5393 ( .A(\RF[30][24] ), .B(n10762), .Y(n193) );
  INVX1 U5394 ( .A(n193), .Y(n4753) );
  AND2X1 U5395 ( .A(\RF[31][58] ), .B(n10764), .Y(n155) );
  INVX1 U5396 ( .A(n155), .Y(n4754) );
  AND2X1 U5397 ( .A(\RF[31][48] ), .B(n10764), .Y(n135) );
  INVX1 U5398 ( .A(n135), .Y(n4755) );
  AND2X1 U5399 ( .A(\RF[0][47] ), .B(n10701), .Y(n2177) );
  INVX1 U5400 ( .A(n2177), .Y(n4756) );
  AND2X1 U5401 ( .A(\RF[0][25] ), .B(n10702), .Y(n2155) );
  INVX1 U5402 ( .A(n2155), .Y(n4757) );
  AND2X1 U5403 ( .A(\RF[0][20] ), .B(n10702), .Y(n2150) );
  INVX1 U5404 ( .A(n2150), .Y(n4758) );
  AND2X1 U5405 ( .A(\RF[0][8] ), .B(n10702), .Y(n2138) );
  INVX1 U5406 ( .A(n2138), .Y(n4759) );
  AND2X1 U5407 ( .A(\RF[1][43] ), .B(n10703), .Y(n2108) );
  INVX1 U5408 ( .A(n2108), .Y(n4760) );
  AND2X1 U5409 ( .A(\RF[1][31] ), .B(n10704), .Y(n2096) );
  INVX1 U5410 ( .A(n2096), .Y(n4761) );
  AND2X1 U5411 ( .A(\RF[1][19] ), .B(n10704), .Y(n2084) );
  INVX1 U5412 ( .A(n2084), .Y(n4762) );
  AND2X1 U5413 ( .A(\RF[1][7] ), .B(n10704), .Y(n2072) );
  INVX1 U5414 ( .A(n2072), .Y(n4763) );
  AND2X1 U5415 ( .A(\RF[2][38] ), .B(n10706), .Y(n2038) );
  INVX1 U5416 ( .A(n2038), .Y(n4764) );
  AND2X1 U5417 ( .A(\RF[2][30] ), .B(n10705), .Y(n2030) );
  INVX1 U5418 ( .A(n2030), .Y(n4765) );
  AND2X1 U5419 ( .A(\RF[2][18] ), .B(n10705), .Y(n2018) );
  INVX1 U5420 ( .A(n2018), .Y(n4766) );
  AND2X1 U5421 ( .A(\RF[2][6] ), .B(n10706), .Y(n2006) );
  INVX1 U5422 ( .A(n2006), .Y(n4767) );
  AND2X1 U5423 ( .A(\RF[3][41] ), .B(n10707), .Y(n1976) );
  INVX1 U5424 ( .A(n1976), .Y(n4768) );
  AND2X1 U5425 ( .A(\RF[3][29] ), .B(n10708), .Y(n1964) );
  INVX1 U5426 ( .A(n1964), .Y(n4769) );
  AND2X1 U5427 ( .A(\RF[3][17] ), .B(n10708), .Y(n1952) );
  INVX1 U5428 ( .A(n1952), .Y(n4770) );
  AND2X1 U5429 ( .A(\RF[3][5] ), .B(n10708), .Y(n1940) );
  INVX1 U5430 ( .A(n1940), .Y(n4771) );
  AND2X1 U5431 ( .A(\RF[4][59] ), .B(n10710), .Y(n1929) );
  INVX1 U5432 ( .A(n1929), .Y(n4772) );
  AND2X1 U5433 ( .A(\RF[4][42] ), .B(n10710), .Y(n1912) );
  INVX1 U5434 ( .A(n1912), .Y(n4773) );
  AND2X1 U5435 ( .A(\RF[4][36] ), .B(n10710), .Y(n1906) );
  INVX1 U5436 ( .A(n1906), .Y(n4774) );
  AND2X1 U5437 ( .A(\RF[4][12] ), .B(n10710), .Y(n1882) );
  INVX1 U5438 ( .A(n1882), .Y(n4775) );
  AND2X1 U5439 ( .A(\RF[5][56] ), .B(n10712), .Y(n1861) );
  INVX1 U5440 ( .A(n1861), .Y(n4776) );
  AND2X1 U5441 ( .A(\RF[5][35] ), .B(n10712), .Y(n1840) );
  INVX1 U5442 ( .A(n1840), .Y(n4777) );
  AND2X1 U5443 ( .A(\RF[5][23] ), .B(n10712), .Y(n1828) );
  INVX1 U5444 ( .A(n1828), .Y(n4778) );
  AND2X1 U5445 ( .A(\RF[5][11] ), .B(n10711), .Y(n1816) );
  INVX1 U5446 ( .A(n1816), .Y(n4779) );
  AND2X1 U5447 ( .A(\RF[6][63] ), .B(n10714), .Y(n1803) );
  INVX1 U5448 ( .A(n1803), .Y(n4780) );
  AND2X1 U5449 ( .A(\RF[6][34] ), .B(n10714), .Y(n1774) );
  INVX1 U5450 ( .A(n1774), .Y(n4781) );
  AND2X1 U5451 ( .A(\RF[6][22] ), .B(n10713), .Y(n1762) );
  INVX1 U5452 ( .A(n1762), .Y(n4782) );
  AND2X1 U5453 ( .A(\RF[6][10] ), .B(n10714), .Y(n1750) );
  INVX1 U5454 ( .A(n1750), .Y(n4783) );
  AND2X1 U5455 ( .A(\RF[7][44] ), .B(n10715), .Y(n1718) );
  INVX1 U5456 ( .A(n1718), .Y(n4784) );
  AND2X1 U5457 ( .A(\RF[7][33] ), .B(n10716), .Y(n1707) );
  INVX1 U5458 ( .A(n1707), .Y(n4785) );
  AND2X1 U5459 ( .A(\RF[7][21] ), .B(n10716), .Y(n1695) );
  INVX1 U5460 ( .A(n1695), .Y(n4786) );
  AND2X1 U5461 ( .A(\RF[7][9] ), .B(n10716), .Y(n1683) );
  INVX1 U5462 ( .A(n1683), .Y(n4787) );
  AND2X1 U5463 ( .A(\RF[8][50] ), .B(n10718), .Y(n1659) );
  INVX1 U5464 ( .A(n1659), .Y(n4788) );
  AND2X1 U5465 ( .A(\RF[9][61] ), .B(n10719), .Y(n1605) );
  INVX1 U5466 ( .A(n1605), .Y(n4789) );
  AND2X1 U5467 ( .A(\RF[9][53] ), .B(n10720), .Y(n1597) );
  INVX1 U5468 ( .A(n1597), .Y(n4790) );
  AND2X1 U5469 ( .A(\RF[9][49] ), .B(n10720), .Y(n1593) );
  INVX1 U5470 ( .A(n1593), .Y(n4791) );
  AND2X1 U5471 ( .A(\RF[10][58] ), .B(n10721), .Y(n1537) );
  INVX1 U5472 ( .A(n1537), .Y(n4792) );
  AND2X1 U5473 ( .A(\RF[10][48] ), .B(n10722), .Y(n1527) );
  INVX1 U5474 ( .A(n1527), .Y(n4793) );
  AND2X1 U5475 ( .A(\RF[11][57] ), .B(n10723), .Y(n1471) );
  INVX1 U5476 ( .A(n1471), .Y(n4794) );
  AND2X1 U5477 ( .A(\RF[11][46] ), .B(n10724), .Y(n1460) );
  INVX1 U5478 ( .A(n1460), .Y(n4795) );
  AND2X1 U5479 ( .A(\RF[11][24] ), .B(n10724), .Y(n1438) );
  INVX1 U5480 ( .A(n1438), .Y(n4796) );
  AND2X1 U5481 ( .A(\RF[12][47] ), .B(n10725), .Y(n1396) );
  INVX1 U5482 ( .A(n1396), .Y(n4797) );
  AND2X1 U5483 ( .A(\RF[12][25] ), .B(n10726), .Y(n1374) );
  INVX1 U5484 ( .A(n1374), .Y(n4798) );
  AND2X1 U5485 ( .A(\RF[12][20] ), .B(n10726), .Y(n1369) );
  INVX1 U5486 ( .A(n1369), .Y(n4799) );
  AND2X1 U5487 ( .A(\RF[12][8] ), .B(n10726), .Y(n1357) );
  INVX1 U5488 ( .A(n1357), .Y(n4800) );
  AND2X1 U5489 ( .A(\RF[13][43] ), .B(n10727), .Y(n1327) );
  INVX1 U5490 ( .A(n1327), .Y(n4801) );
  AND2X1 U5491 ( .A(\RF[13][31] ), .B(n10728), .Y(n1315) );
  INVX1 U5492 ( .A(n1315), .Y(n4802) );
  AND2X1 U5493 ( .A(\RF[13][19] ), .B(n10728), .Y(n1303) );
  INVX1 U5494 ( .A(n1303), .Y(n4803) );
  AND2X1 U5495 ( .A(\RF[13][7] ), .B(n10728), .Y(n1291) );
  INVX1 U5496 ( .A(n1291), .Y(n4804) );
  AND2X1 U5497 ( .A(\RF[14][38] ), .B(n10730), .Y(n1257) );
  INVX1 U5498 ( .A(n1257), .Y(n4805) );
  AND2X1 U5499 ( .A(\RF[14][30] ), .B(n10729), .Y(n1249) );
  INVX1 U5500 ( .A(n1249), .Y(n4806) );
  AND2X1 U5501 ( .A(\RF[14][18] ), .B(n10729), .Y(n1237) );
  INVX1 U5502 ( .A(n1237), .Y(n4807) );
  AND2X1 U5503 ( .A(\RF[14][6] ), .B(n10730), .Y(n1225) );
  INVX1 U5504 ( .A(n1225), .Y(n4808) );
  AND2X1 U5505 ( .A(\RF[15][41] ), .B(n10731), .Y(n1194) );
  INVX1 U5506 ( .A(n1194), .Y(n4809) );
  AND2X1 U5507 ( .A(\RF[15][29] ), .B(n10732), .Y(n1182) );
  INVX1 U5508 ( .A(n1182), .Y(n4810) );
  AND2X1 U5509 ( .A(\RF[15][17] ), .B(n10732), .Y(n1170) );
  INVX1 U5510 ( .A(n1170), .Y(n4811) );
  AND2X1 U5511 ( .A(\RF[15][5] ), .B(n10732), .Y(n1158) );
  INVX1 U5512 ( .A(n1158), .Y(n4812) );
  AND2X1 U5513 ( .A(\RF[16][59] ), .B(n10734), .Y(n1147) );
  INVX1 U5514 ( .A(n1147), .Y(n4813) );
  AND2X1 U5515 ( .A(\RF[16][42] ), .B(n10734), .Y(n1130) );
  INVX1 U5516 ( .A(n1130), .Y(n4814) );
  AND2X1 U5517 ( .A(\RF[16][36] ), .B(n10734), .Y(n1124) );
  INVX1 U5518 ( .A(n1124), .Y(n4815) );
  AND2X1 U5519 ( .A(\RF[16][12] ), .B(n10734), .Y(n1100) );
  INVX1 U5520 ( .A(n1100), .Y(n4816) );
  AND2X1 U5521 ( .A(\RF[17][56] ), .B(n10736), .Y(n1079) );
  INVX1 U5522 ( .A(n1079), .Y(n4817) );
  AND2X1 U5523 ( .A(\RF[17][35] ), .B(n10736), .Y(n1058) );
  INVX1 U5524 ( .A(n1058), .Y(n4818) );
  AND2X1 U5525 ( .A(\RF[17][23] ), .B(n10736), .Y(n1046) );
  INVX1 U5526 ( .A(n1046), .Y(n4819) );
  AND2X1 U5527 ( .A(\RF[17][11] ), .B(n10735), .Y(n1034) );
  INVX1 U5528 ( .A(n1034), .Y(n4820) );
  AND2X1 U5529 ( .A(\RF[18][63] ), .B(n10738), .Y(n1021) );
  INVX1 U5530 ( .A(n1021), .Y(n4821) );
  AND2X1 U5531 ( .A(\RF[18][34] ), .B(n10738), .Y(n992) );
  INVX1 U5532 ( .A(n992), .Y(n4822) );
  AND2X1 U5533 ( .A(\RF[18][22] ), .B(n10737), .Y(n980) );
  INVX1 U5534 ( .A(n980), .Y(n4823) );
  AND2X1 U5535 ( .A(\RF[18][10] ), .B(n10738), .Y(n968) );
  INVX1 U5536 ( .A(n968), .Y(n4824) );
  AND2X1 U5537 ( .A(\RF[19][44] ), .B(n10739), .Y(n937) );
  INVX1 U5538 ( .A(n937), .Y(n4825) );
  AND2X1 U5539 ( .A(\RF[19][33] ), .B(n10740), .Y(n926) );
  INVX1 U5540 ( .A(n926), .Y(n4826) );
  AND2X1 U5541 ( .A(\RF[19][21] ), .B(n10740), .Y(n914) );
  INVX1 U5542 ( .A(n914), .Y(n4827) );
  AND2X1 U5543 ( .A(\RF[19][9] ), .B(n10740), .Y(n902) );
  INVX1 U5544 ( .A(n902), .Y(n4828) );
  AND2X1 U5545 ( .A(\RF[20][50] ), .B(n10742), .Y(n878) );
  INVX1 U5546 ( .A(n878), .Y(n4829) );
  AND2X1 U5547 ( .A(\RF[21][61] ), .B(n10743), .Y(n824) );
  INVX1 U5548 ( .A(n824), .Y(n4830) );
  AND2X1 U5549 ( .A(\RF[21][53] ), .B(n10744), .Y(n816) );
  INVX1 U5550 ( .A(n816), .Y(n4831) );
  AND2X1 U5551 ( .A(\RF[21][49] ), .B(n10744), .Y(n812) );
  INVX1 U5552 ( .A(n812), .Y(n4832) );
  AND2X1 U5553 ( .A(\RF[22][58] ), .B(n10745), .Y(n756) );
  INVX1 U5554 ( .A(n756), .Y(n4833) );
  AND2X1 U5555 ( .A(\RF[22][48] ), .B(n10746), .Y(n746) );
  INVX1 U5556 ( .A(n746), .Y(n4834) );
  AND2X1 U5557 ( .A(\RF[23][57] ), .B(n10747), .Y(n689) );
  INVX1 U5558 ( .A(n689), .Y(n4835) );
  AND2X1 U5559 ( .A(\RF[23][46] ), .B(n10748), .Y(n678) );
  INVX1 U5560 ( .A(n678), .Y(n4836) );
  AND2X1 U5561 ( .A(\RF[23][24] ), .B(n10748), .Y(n656) );
  INVX1 U5562 ( .A(n656), .Y(n4837) );
  AND2X1 U5563 ( .A(\RF[24][59] ), .B(n10750), .Y(n624) );
  INVX1 U5564 ( .A(n624), .Y(n4838) );
  AND2X1 U5565 ( .A(\RF[24][42] ), .B(n10750), .Y(n607) );
  INVX1 U5566 ( .A(n607), .Y(n4839) );
  AND2X1 U5567 ( .A(\RF[24][36] ), .B(n10750), .Y(n601) );
  INVX1 U5568 ( .A(n601), .Y(n4840) );
  AND2X1 U5569 ( .A(\RF[24][12] ), .B(n10750), .Y(n577) );
  INVX1 U5570 ( .A(n577), .Y(n4841) );
  AND2X1 U5571 ( .A(\RF[25][56] ), .B(n10752), .Y(n555) );
  INVX1 U5572 ( .A(n555), .Y(n4842) );
  AND2X1 U5573 ( .A(\RF[25][35] ), .B(n10752), .Y(n534) );
  INVX1 U5574 ( .A(n534), .Y(n4843) );
  AND2X1 U5575 ( .A(\RF[25][23] ), .B(n10752), .Y(n522) );
  INVX1 U5576 ( .A(n522), .Y(n4844) );
  AND2X1 U5577 ( .A(\RF[25][11] ), .B(n10751), .Y(n510) );
  INVX1 U5578 ( .A(n510), .Y(n4845) );
  AND2X1 U5579 ( .A(\RF[26][63] ), .B(n10754), .Y(n496) );
  INVX1 U5580 ( .A(n496), .Y(n4846) );
  AND2X1 U5581 ( .A(\RF[26][34] ), .B(n10754), .Y(n467) );
  INVX1 U5582 ( .A(n467), .Y(n4847) );
  AND2X1 U5583 ( .A(\RF[26][22] ), .B(n10753), .Y(n455) );
  INVX1 U5584 ( .A(n455), .Y(n4848) );
  AND2X1 U5585 ( .A(\RF[26][10] ), .B(n10754), .Y(n443) );
  INVX1 U5586 ( .A(n443), .Y(n4849) );
  AND2X1 U5587 ( .A(\RF[27][44] ), .B(n10755), .Y(n411) );
  INVX1 U5588 ( .A(n411), .Y(n4850) );
  AND2X1 U5589 ( .A(\RF[27][33] ), .B(n10756), .Y(n400) );
  INVX1 U5590 ( .A(n400), .Y(n4851) );
  AND2X1 U5591 ( .A(\RF[27][21] ), .B(n10756), .Y(n388) );
  INVX1 U5592 ( .A(n388), .Y(n4852) );
  AND2X1 U5593 ( .A(\RF[27][9] ), .B(n10756), .Y(n376) );
  INVX1 U5594 ( .A(n376), .Y(n4853) );
  AND2X1 U5595 ( .A(\RF[28][50] ), .B(n10758), .Y(n351) );
  INVX1 U5596 ( .A(n351), .Y(n4854) );
  AND2X1 U5597 ( .A(\RF[29][61] ), .B(n10759), .Y(n296) );
  INVX1 U5598 ( .A(n296), .Y(n4855) );
  AND2X1 U5599 ( .A(\RF[29][53] ), .B(n10760), .Y(n288) );
  INVX1 U5600 ( .A(n288), .Y(n4856) );
  AND2X1 U5601 ( .A(\RF[29][49] ), .B(n10760), .Y(n284) );
  INVX1 U5602 ( .A(n284), .Y(n4857) );
  AND2X1 U5603 ( .A(\RF[30][58] ), .B(n10761), .Y(n227) );
  INVX1 U5604 ( .A(n227), .Y(n4858) );
  AND2X1 U5605 ( .A(\RF[30][48] ), .B(n10762), .Y(n217) );
  INVX1 U5606 ( .A(n217), .Y(n4859) );
  AND2X1 U5607 ( .A(\RF[31][57] ), .B(n10763), .Y(n153) );
  INVX1 U5608 ( .A(n153), .Y(n4860) );
  AND2X1 U5609 ( .A(\RF[31][46] ), .B(n10764), .Y(n131) );
  INVX1 U5610 ( .A(n131), .Y(n4861) );
  AND2X1 U5611 ( .A(\RF[31][24] ), .B(n10764), .Y(n87) );
  INVX1 U5612 ( .A(n87), .Y(n4862) );
  AND2X1 U5613 ( .A(\RF[0][45] ), .B(n10701), .Y(n2175) );
  INVX1 U5614 ( .A(n2175), .Y(n4863) );
  AND2X1 U5615 ( .A(\RF[0][32] ), .B(n10702), .Y(n2162) );
  INVX1 U5616 ( .A(n2162), .Y(n4864) );
  AND2X1 U5617 ( .A(\RF[0][13] ), .B(n10702), .Y(n2143) );
  INVX1 U5618 ( .A(n2143), .Y(n4865) );
  AND2X1 U5619 ( .A(\RF[0][1] ), .B(n10702), .Y(n2131) );
  INVX1 U5620 ( .A(n2131), .Y(n4866) );
  AND2X1 U5621 ( .A(\RF[0][0] ), .B(n10702), .Y(n2130) );
  INVX1 U5622 ( .A(n2130), .Y(n4867) );
  AND2X1 U5623 ( .A(\RF[1][37] ), .B(n10704), .Y(n2102) );
  INVX1 U5624 ( .A(n2102), .Y(n4868) );
  AND2X1 U5625 ( .A(\RF[1][26] ), .B(n10703), .Y(n2091) );
  INVX1 U5626 ( .A(n2091), .Y(n4869) );
  AND2X1 U5627 ( .A(\RF[1][14] ), .B(n10704), .Y(n2079) );
  INVX1 U5628 ( .A(n2079), .Y(n4870) );
  AND2X1 U5629 ( .A(\RF[1][2] ), .B(n10704), .Y(n2067) );
  INVX1 U5630 ( .A(n2067), .Y(n4871) );
  AND2X1 U5631 ( .A(\RF[2][39] ), .B(n10706), .Y(n2039) );
  INVX1 U5632 ( .A(n2039), .Y(n4872) );
  AND2X1 U5633 ( .A(\RF[2][27] ), .B(n10706), .Y(n2027) );
  INVX1 U5634 ( .A(n2027), .Y(n4873) );
  AND2X1 U5635 ( .A(\RF[2][15] ), .B(n10706), .Y(n2015) );
  INVX1 U5636 ( .A(n2015), .Y(n4874) );
  AND2X1 U5637 ( .A(\RF[2][3] ), .B(n10706), .Y(n2003) );
  INVX1 U5638 ( .A(n2003), .Y(n4875) );
  AND2X1 U5639 ( .A(\RF[3][40] ), .B(n10708), .Y(n1975) );
  INVX1 U5640 ( .A(n1975), .Y(n4876) );
  AND2X1 U5641 ( .A(\RF[3][28] ), .B(n10707), .Y(n1963) );
  INVX1 U5642 ( .A(n1963), .Y(n4877) );
  AND2X1 U5643 ( .A(\RF[3][16] ), .B(n10708), .Y(n1951) );
  INVX1 U5644 ( .A(n1951), .Y(n4878) );
  AND2X1 U5645 ( .A(\RF[3][4] ), .B(n10708), .Y(n1939) );
  INVX1 U5646 ( .A(n1939), .Y(n4879) );
  AND2X1 U5647 ( .A(\RF[4][57] ), .B(n10710), .Y(n1927) );
  INVX1 U5648 ( .A(n1927), .Y(n4880) );
  AND2X1 U5649 ( .A(\RF[4][46] ), .B(n10709), .Y(n1916) );
  INVX1 U5650 ( .A(n1916), .Y(n4881) );
  AND2X1 U5651 ( .A(\RF[4][24] ), .B(n10710), .Y(n1894) );
  INVX1 U5652 ( .A(n1894), .Y(n4882) );
  AND2X1 U5653 ( .A(\RF[5][58] ), .B(n10712), .Y(n1863) );
  INVX1 U5654 ( .A(n1863), .Y(n4883) );
  AND2X1 U5655 ( .A(\RF[5][48] ), .B(n10712), .Y(n1853) );
  INVX1 U5656 ( .A(n1853), .Y(n4884) );
  AND2X1 U5657 ( .A(\RF[6][61] ), .B(n10714), .Y(n1801) );
  INVX1 U5658 ( .A(n1801), .Y(n4885) );
  AND2X1 U5659 ( .A(\RF[6][53] ), .B(n10714), .Y(n1793) );
  INVX1 U5660 ( .A(n1793), .Y(n4886) );
  AND2X1 U5661 ( .A(\RF[6][49] ), .B(n10714), .Y(n1789) );
  INVX1 U5662 ( .A(n1789), .Y(n4887) );
  AND2X1 U5663 ( .A(\RF[7][50] ), .B(n10716), .Y(n1724) );
  INVX1 U5664 ( .A(n1724), .Y(n4888) );
  AND2X1 U5665 ( .A(\RF[8][44] ), .B(n10717), .Y(n1653) );
  INVX1 U5666 ( .A(n1653), .Y(n4889) );
  AND2X1 U5667 ( .A(\RF[8][33] ), .B(n10718), .Y(n1642) );
  INVX1 U5668 ( .A(n1642), .Y(n4890) );
  AND2X1 U5669 ( .A(\RF[8][21] ), .B(n10718), .Y(n1630) );
  INVX1 U5670 ( .A(n1630), .Y(n4891) );
  AND2X1 U5671 ( .A(\RF[8][9] ), .B(n10718), .Y(n1618) );
  INVX1 U5672 ( .A(n1618), .Y(n4892) );
  AND2X1 U5673 ( .A(\RF[9][63] ), .B(n10720), .Y(n1607) );
  INVX1 U5674 ( .A(n1607), .Y(n4893) );
  AND2X1 U5675 ( .A(\RF[9][34] ), .B(n10720), .Y(n1578) );
  INVX1 U5676 ( .A(n1578), .Y(n4894) );
  AND2X1 U5677 ( .A(\RF[9][22] ), .B(n10719), .Y(n1566) );
  INVX1 U5678 ( .A(n1566), .Y(n4895) );
  AND2X1 U5679 ( .A(\RF[9][10] ), .B(n10720), .Y(n1554) );
  INVX1 U5680 ( .A(n1554), .Y(n4896) );
  AND2X1 U5681 ( .A(\RF[10][56] ), .B(n10722), .Y(n1535) );
  INVX1 U5682 ( .A(n1535), .Y(n4897) );
  AND2X1 U5683 ( .A(\RF[10][35] ), .B(n10722), .Y(n1514) );
  INVX1 U5684 ( .A(n1514), .Y(n4898) );
  AND2X1 U5685 ( .A(\RF[10][23] ), .B(n10722), .Y(n1502) );
  INVX1 U5686 ( .A(n1502), .Y(n4899) );
  AND2X1 U5687 ( .A(\RF[10][11] ), .B(n10721), .Y(n1490) );
  INVX1 U5688 ( .A(n1490), .Y(n4900) );
  AND2X1 U5689 ( .A(\RF[11][59] ), .B(n10724), .Y(n1473) );
  INVX1 U5690 ( .A(n1473), .Y(n4901) );
  AND2X1 U5691 ( .A(\RF[11][42] ), .B(n10724), .Y(n1456) );
  INVX1 U5692 ( .A(n1456), .Y(n4902) );
  AND2X1 U5693 ( .A(\RF[11][36] ), .B(n10724), .Y(n1450) );
  INVX1 U5694 ( .A(n1450), .Y(n4903) );
  AND2X1 U5695 ( .A(\RF[11][12] ), .B(n10723), .Y(n1426) );
  INVX1 U5696 ( .A(n1426), .Y(n4904) );
  AND2X1 U5697 ( .A(\RF[12][45] ), .B(n10725), .Y(n1394) );
  INVX1 U5698 ( .A(n1394), .Y(n4905) );
  AND2X1 U5699 ( .A(\RF[12][32] ), .B(n10726), .Y(n1381) );
  INVX1 U5700 ( .A(n1381), .Y(n4906) );
  AND2X1 U5701 ( .A(\RF[12][13] ), .B(n10726), .Y(n1362) );
  INVX1 U5702 ( .A(n1362), .Y(n4907) );
  AND2X1 U5703 ( .A(\RF[12][1] ), .B(n10726), .Y(n1350) );
  INVX1 U5704 ( .A(n1350), .Y(n4908) );
  AND2X1 U5705 ( .A(\RF[12][0] ), .B(n10726), .Y(n1349) );
  INVX1 U5706 ( .A(n1349), .Y(n4909) );
  AND2X1 U5707 ( .A(\RF[13][37] ), .B(n10728), .Y(n1321) );
  INVX1 U5708 ( .A(n1321), .Y(n4910) );
  AND2X1 U5709 ( .A(\RF[13][26] ), .B(n10727), .Y(n1310) );
  INVX1 U5710 ( .A(n1310), .Y(n4911) );
  AND2X1 U5711 ( .A(\RF[13][14] ), .B(n10728), .Y(n1298) );
  INVX1 U5712 ( .A(n1298), .Y(n4912) );
  AND2X1 U5713 ( .A(\RF[13][2] ), .B(n10728), .Y(n1286) );
  INVX1 U5714 ( .A(n1286), .Y(n4913) );
  AND2X1 U5715 ( .A(\RF[14][39] ), .B(n10730), .Y(n1258) );
  INVX1 U5716 ( .A(n1258), .Y(n4914) );
  AND2X1 U5717 ( .A(\RF[14][27] ), .B(n10730), .Y(n1246) );
  INVX1 U5718 ( .A(n1246), .Y(n4915) );
  AND2X1 U5719 ( .A(\RF[14][15] ), .B(n10730), .Y(n1234) );
  INVX1 U5720 ( .A(n1234), .Y(n4916) );
  AND2X1 U5721 ( .A(\RF[14][3] ), .B(n10730), .Y(n1222) );
  INVX1 U5722 ( .A(n1222), .Y(n4917) );
  AND2X1 U5723 ( .A(\RF[15][40] ), .B(n10732), .Y(n1193) );
  INVX1 U5724 ( .A(n1193), .Y(n4918) );
  AND2X1 U5725 ( .A(\RF[15][28] ), .B(n10731), .Y(n1181) );
  INVX1 U5726 ( .A(n1181), .Y(n4919) );
  AND2X1 U5727 ( .A(\RF[15][16] ), .B(n10732), .Y(n1169) );
  INVX1 U5728 ( .A(n1169), .Y(n4920) );
  AND2X1 U5729 ( .A(\RF[15][4] ), .B(n10732), .Y(n1157) );
  INVX1 U5730 ( .A(n1157), .Y(n4921) );
  AND2X1 U5731 ( .A(\RF[16][57] ), .B(n10734), .Y(n1145) );
  INVX1 U5732 ( .A(n1145), .Y(n4922) );
  AND2X1 U5733 ( .A(\RF[16][46] ), .B(n10733), .Y(n1134) );
  INVX1 U5734 ( .A(n1134), .Y(n4923) );
  AND2X1 U5735 ( .A(\RF[16][24] ), .B(n10734), .Y(n1112) );
  INVX1 U5736 ( .A(n1112), .Y(n4924) );
  AND2X1 U5737 ( .A(\RF[17][58] ), .B(n10736), .Y(n1081) );
  INVX1 U5738 ( .A(n1081), .Y(n4925) );
  AND2X1 U5739 ( .A(\RF[17][48] ), .B(n10736), .Y(n1071) );
  INVX1 U5740 ( .A(n1071), .Y(n4926) );
  AND2X1 U5741 ( .A(\RF[18][61] ), .B(n10738), .Y(n1019) );
  INVX1 U5742 ( .A(n1019), .Y(n4927) );
  AND2X1 U5743 ( .A(\RF[18][53] ), .B(n10738), .Y(n1011) );
  INVX1 U5744 ( .A(n1011), .Y(n4928) );
  AND2X1 U5745 ( .A(\RF[18][49] ), .B(n10738), .Y(n1007) );
  INVX1 U5746 ( .A(n1007), .Y(n4929) );
  AND2X1 U5747 ( .A(\RF[19][50] ), .B(n10740), .Y(n943) );
  INVX1 U5748 ( .A(n943), .Y(n4930) );
  AND2X1 U5749 ( .A(\RF[20][44] ), .B(n10741), .Y(n872) );
  INVX1 U5750 ( .A(n872), .Y(n4931) );
  AND2X1 U5751 ( .A(\RF[20][33] ), .B(n10742), .Y(n861) );
  INVX1 U5752 ( .A(n861), .Y(n4932) );
  AND2X1 U5753 ( .A(\RF[20][21] ), .B(n10742), .Y(n849) );
  INVX1 U5754 ( .A(n849), .Y(n4933) );
  AND2X1 U5755 ( .A(\RF[20][9] ), .B(n10742), .Y(n837) );
  INVX1 U5756 ( .A(n837), .Y(n4934) );
  AND2X1 U5757 ( .A(\RF[21][63] ), .B(n10744), .Y(n826) );
  INVX1 U5758 ( .A(n826), .Y(n4935) );
  AND2X1 U5759 ( .A(\RF[21][34] ), .B(n10744), .Y(n797) );
  INVX1 U5760 ( .A(n797), .Y(n4936) );
  AND2X1 U5761 ( .A(\RF[21][22] ), .B(n10743), .Y(n785) );
  INVX1 U5762 ( .A(n785), .Y(n4937) );
  AND2X1 U5763 ( .A(\RF[21][10] ), .B(n10744), .Y(n773) );
  INVX1 U5764 ( .A(n773), .Y(n4938) );
  AND2X1 U5765 ( .A(\RF[22][56] ), .B(n10746), .Y(n754) );
  INVX1 U5766 ( .A(n754), .Y(n4939) );
  AND2X1 U5767 ( .A(\RF[22][35] ), .B(n10746), .Y(n733) );
  INVX1 U5768 ( .A(n733), .Y(n4940) );
  AND2X1 U5769 ( .A(\RF[22][23] ), .B(n10746), .Y(n721) );
  INVX1 U5770 ( .A(n721), .Y(n4941) );
  AND2X1 U5771 ( .A(\RF[22][11] ), .B(n10745), .Y(n709) );
  INVX1 U5772 ( .A(n709), .Y(n4942) );
  AND2X1 U5773 ( .A(\RF[23][59] ), .B(n10748), .Y(n691) );
  INVX1 U5774 ( .A(n691), .Y(n4943) );
  AND2X1 U5775 ( .A(\RF[23][42] ), .B(n10748), .Y(n674) );
  INVX1 U5776 ( .A(n674), .Y(n4944) );
  AND2X1 U5777 ( .A(\RF[23][36] ), .B(n10748), .Y(n668) );
  INVX1 U5778 ( .A(n668), .Y(n4945) );
  AND2X1 U5779 ( .A(\RF[23][12] ), .B(n10747), .Y(n644) );
  INVX1 U5780 ( .A(n644), .Y(n4946) );
  AND2X1 U5781 ( .A(\RF[24][57] ), .B(n10750), .Y(n622) );
  INVX1 U5782 ( .A(n622), .Y(n4947) );
  AND2X1 U5783 ( .A(\RF[24][46] ), .B(n10749), .Y(n611) );
  INVX1 U5784 ( .A(n611), .Y(n4948) );
  AND2X1 U5785 ( .A(\RF[24][24] ), .B(n10750), .Y(n589) );
  INVX1 U5786 ( .A(n589), .Y(n4949) );
  AND2X1 U5787 ( .A(\RF[25][58] ), .B(n10752), .Y(n557) );
  INVX1 U5788 ( .A(n557), .Y(n4950) );
  AND2X1 U5789 ( .A(\RF[25][48] ), .B(n10752), .Y(n547) );
  INVX1 U5790 ( .A(n547), .Y(n4951) );
  AND2X1 U5791 ( .A(\RF[26][61] ), .B(n10754), .Y(n494) );
  INVX1 U5792 ( .A(n494), .Y(n4952) );
  AND2X1 U5793 ( .A(\RF[26][53] ), .B(n10754), .Y(n486) );
  INVX1 U5794 ( .A(n486), .Y(n4953) );
  AND2X1 U5795 ( .A(\RF[26][49] ), .B(n10754), .Y(n482) );
  INVX1 U5796 ( .A(n482), .Y(n4954) );
  AND2X1 U5797 ( .A(\RF[27][50] ), .B(n10756), .Y(n417) );
  INVX1 U5798 ( .A(n417), .Y(n4955) );
  AND2X1 U5799 ( .A(\RF[28][44] ), .B(n10757), .Y(n345) );
  INVX1 U5800 ( .A(n345), .Y(n4956) );
  AND2X1 U5801 ( .A(\RF[28][33] ), .B(n10758), .Y(n334) );
  INVX1 U5802 ( .A(n334), .Y(n4957) );
  AND2X1 U5803 ( .A(\RF[28][21] ), .B(n10758), .Y(n322) );
  INVX1 U5804 ( .A(n322), .Y(n4958) );
  AND2X1 U5805 ( .A(\RF[28][9] ), .B(n10758), .Y(n310) );
  INVX1 U5806 ( .A(n310), .Y(n4959) );
  AND2X1 U5807 ( .A(\RF[29][63] ), .B(n10760), .Y(n298) );
  INVX1 U5808 ( .A(n298), .Y(n4960) );
  AND2X1 U5809 ( .A(\RF[29][34] ), .B(n10760), .Y(n269) );
  INVX1 U5810 ( .A(n269), .Y(n4961) );
  AND2X1 U5811 ( .A(\RF[29][22] ), .B(n10759), .Y(n257) );
  INVX1 U5812 ( .A(n257), .Y(n4962) );
  AND2X1 U5813 ( .A(\RF[29][10] ), .B(n10760), .Y(n245) );
  INVX1 U5814 ( .A(n245), .Y(n4963) );
  AND2X1 U5815 ( .A(\RF[30][56] ), .B(n10762), .Y(n225) );
  INVX1 U5816 ( .A(n225), .Y(n4964) );
  AND2X1 U5817 ( .A(\RF[30][35] ), .B(n10762), .Y(n204) );
  INVX1 U5818 ( .A(n204), .Y(n4965) );
  AND2X1 U5819 ( .A(\RF[30][23] ), .B(n10762), .Y(n192) );
  INVX1 U5820 ( .A(n192), .Y(n4966) );
  AND2X1 U5821 ( .A(\RF[30][11] ), .B(n10761), .Y(n180) );
  INVX1 U5822 ( .A(n180), .Y(n4967) );
  AND2X1 U5823 ( .A(\RF[31][59] ), .B(n10764), .Y(n157) );
  INVX1 U5824 ( .A(n157), .Y(n4968) );
  AND2X1 U5825 ( .A(\RF[31][42] ), .B(n10764), .Y(n123) );
  INVX1 U5826 ( .A(n123), .Y(n4969) );
  AND2X1 U5827 ( .A(\RF[31][36] ), .B(n10764), .Y(n111) );
  INVX1 U5828 ( .A(n111), .Y(n4970) );
  AND2X1 U5829 ( .A(\RF[31][12] ), .B(n10763), .Y(n63) );
  INVX1 U5830 ( .A(n63), .Y(n4971) );
  AND2X1 U5831 ( .A(\RF[0][37] ), .B(n10701), .Y(n2167) );
  INVX1 U5832 ( .A(n2167), .Y(n4972) );
  AND2X1 U5833 ( .A(\RF[0][26] ), .B(n10701), .Y(n2156) );
  INVX1 U5834 ( .A(n2156), .Y(n4973) );
  AND2X1 U5835 ( .A(\RF[0][14] ), .B(n10702), .Y(n2144) );
  INVX1 U5836 ( .A(n2144), .Y(n4974) );
  AND2X1 U5837 ( .A(\RF[0][2] ), .B(n10702), .Y(n2132) );
  INVX1 U5838 ( .A(n2132), .Y(n4975) );
  AND2X1 U5839 ( .A(\RF[1][45] ), .B(n10703), .Y(n2110) );
  INVX1 U5840 ( .A(n2110), .Y(n4976) );
  AND2X1 U5841 ( .A(\RF[1][32] ), .B(n10703), .Y(n2097) );
  INVX1 U5842 ( .A(n2097), .Y(n4977) );
  AND2X1 U5843 ( .A(\RF[1][13] ), .B(n10704), .Y(n2078) );
  INVX1 U5844 ( .A(n2078), .Y(n4978) );
  AND2X1 U5845 ( .A(\RF[1][1] ), .B(n10704), .Y(n2066) );
  INVX1 U5846 ( .A(n2066), .Y(n4979) );
  AND2X1 U5847 ( .A(\RF[1][0] ), .B(n10704), .Y(n2065) );
  INVX1 U5848 ( .A(n2065), .Y(n4980) );
  AND2X1 U5849 ( .A(\RF[2][40] ), .B(n10705), .Y(n2040) );
  INVX1 U5850 ( .A(n2040), .Y(n4981) );
  AND2X1 U5851 ( .A(\RF[2][28] ), .B(n10706), .Y(n2028) );
  INVX1 U5852 ( .A(n2028), .Y(n4982) );
  AND2X1 U5853 ( .A(\RF[2][16] ), .B(n10706), .Y(n2016) );
  INVX1 U5854 ( .A(n2016), .Y(n4983) );
  AND2X1 U5855 ( .A(\RF[2][4] ), .B(n10706), .Y(n2004) );
  INVX1 U5856 ( .A(n2004), .Y(n4984) );
  AND2X1 U5857 ( .A(\RF[3][39] ), .B(n10707), .Y(n1974) );
  INVX1 U5858 ( .A(n1974), .Y(n4985) );
  AND2X1 U5859 ( .A(\RF[3][27] ), .B(n10707), .Y(n1962) );
  INVX1 U5860 ( .A(n1962), .Y(n4986) );
  AND2X1 U5861 ( .A(\RF[3][15] ), .B(n10708), .Y(n1950) );
  INVX1 U5862 ( .A(n1950), .Y(n4987) );
  AND2X1 U5863 ( .A(\RF[3][3] ), .B(n10708), .Y(n1938) );
  INVX1 U5864 ( .A(n1938), .Y(n4988) );
  AND2X1 U5865 ( .A(\RF[4][58] ), .B(n10710), .Y(n1928) );
  INVX1 U5866 ( .A(n1928), .Y(n4989) );
  AND2X1 U5867 ( .A(\RF[4][48] ), .B(n10709), .Y(n1918) );
  INVX1 U5868 ( .A(n1918), .Y(n4990) );
  AND2X1 U5869 ( .A(\RF[5][57] ), .B(n10712), .Y(n1862) );
  INVX1 U5870 ( .A(n1862), .Y(n4991) );
  AND2X1 U5871 ( .A(\RF[5][46] ), .B(n10712), .Y(n1851) );
  INVX1 U5872 ( .A(n1851), .Y(n4992) );
  AND2X1 U5873 ( .A(\RF[5][24] ), .B(n10712), .Y(n1829) );
  INVX1 U5874 ( .A(n1829), .Y(n4993) );
  AND2X1 U5875 ( .A(\RF[6][50] ), .B(n10714), .Y(n1790) );
  INVX1 U5876 ( .A(n1790), .Y(n4994) );
  AND2X1 U5877 ( .A(\RF[7][61] ), .B(n10716), .Y(n1735) );
  INVX1 U5878 ( .A(n1735), .Y(n4995) );
  AND2X1 U5879 ( .A(\RF[7][53] ), .B(n10716), .Y(n1727) );
  INVX1 U5880 ( .A(n1727), .Y(n4996) );
  AND2X1 U5881 ( .A(\RF[7][49] ), .B(n10716), .Y(n1723) );
  INVX1 U5882 ( .A(n1723), .Y(n4997) );
  AND2X1 U5883 ( .A(\RF[8][63] ), .B(n10718), .Y(n1672) );
  INVX1 U5884 ( .A(n1672), .Y(n4998) );
  AND2X1 U5885 ( .A(\RF[8][34] ), .B(n10718), .Y(n1643) );
  INVX1 U5886 ( .A(n1643), .Y(n4999) );
  AND2X1 U5887 ( .A(\RF[8][22] ), .B(n10717), .Y(n1631) );
  INVX1 U5888 ( .A(n1631), .Y(n5000) );
  AND2X1 U5889 ( .A(\RF[8][10] ), .B(n10718), .Y(n1619) );
  INVX1 U5890 ( .A(n1619), .Y(n5001) );
  AND2X1 U5891 ( .A(\RF[9][44] ), .B(n10719), .Y(n1588) );
  INVX1 U5892 ( .A(n1588), .Y(n5002) );
  AND2X1 U5893 ( .A(\RF[9][33] ), .B(n10720), .Y(n1577) );
  INVX1 U5894 ( .A(n1577), .Y(n5003) );
  AND2X1 U5895 ( .A(\RF[9][21] ), .B(n10720), .Y(n1565) );
  INVX1 U5896 ( .A(n1565), .Y(n5004) );
  AND2X1 U5897 ( .A(\RF[9][9] ), .B(n10720), .Y(n1553) );
  INVX1 U5898 ( .A(n1553), .Y(n5005) );
  AND2X1 U5899 ( .A(\RF[10][59] ), .B(n10722), .Y(n1538) );
  INVX1 U5900 ( .A(n1538), .Y(n5006) );
  AND2X1 U5901 ( .A(\RF[10][42] ), .B(n10722), .Y(n1521) );
  INVX1 U5902 ( .A(n1521), .Y(n5007) );
  AND2X1 U5903 ( .A(\RF[10][36] ), .B(n10721), .Y(n1515) );
  INVX1 U5904 ( .A(n1515), .Y(n5008) );
  AND2X1 U5905 ( .A(\RF[10][12] ), .B(n10721), .Y(n1491) );
  INVX1 U5906 ( .A(n1491), .Y(n5009) );
  AND2X1 U5907 ( .A(\RF[11][56] ), .B(n10724), .Y(n1470) );
  INVX1 U5908 ( .A(n1470), .Y(n5010) );
  AND2X1 U5909 ( .A(\RF[11][35] ), .B(n10723), .Y(n1449) );
  INVX1 U5910 ( .A(n1449), .Y(n5011) );
  AND2X1 U5911 ( .A(\RF[11][23] ), .B(n10724), .Y(n1437) );
  INVX1 U5912 ( .A(n1437), .Y(n5012) );
  AND2X1 U5913 ( .A(\RF[11][11] ), .B(n10723), .Y(n1425) );
  INVX1 U5914 ( .A(n1425), .Y(n5013) );
  AND2X1 U5915 ( .A(\RF[12][37] ), .B(n10725), .Y(n1386) );
  INVX1 U5916 ( .A(n1386), .Y(n5014) );
  AND2X1 U5917 ( .A(\RF[12][26] ), .B(n10725), .Y(n1375) );
  INVX1 U5918 ( .A(n1375), .Y(n5015) );
  AND2X1 U5919 ( .A(\RF[12][14] ), .B(n10726), .Y(n1363) );
  INVX1 U5920 ( .A(n1363), .Y(n5016) );
  AND2X1 U5921 ( .A(\RF[12][2] ), .B(n10726), .Y(n1351) );
  INVX1 U5922 ( .A(n1351), .Y(n5017) );
  AND2X1 U5923 ( .A(\RF[13][45] ), .B(n10727), .Y(n1329) );
  INVX1 U5924 ( .A(n1329), .Y(n5018) );
  AND2X1 U5925 ( .A(\RF[13][32] ), .B(n10727), .Y(n1316) );
  INVX1 U5926 ( .A(n1316), .Y(n5019) );
  AND2X1 U5927 ( .A(\RF[13][13] ), .B(n10728), .Y(n1297) );
  INVX1 U5928 ( .A(n1297), .Y(n5020) );
  AND2X1 U5929 ( .A(\RF[13][1] ), .B(n10728), .Y(n1285) );
  INVX1 U5930 ( .A(n1285), .Y(n5021) );
  AND2X1 U5931 ( .A(\RF[13][0] ), .B(n10728), .Y(n1284) );
  INVX1 U5932 ( .A(n1284), .Y(n5022) );
  AND2X1 U5933 ( .A(\RF[14][40] ), .B(n10729), .Y(n1259) );
  INVX1 U5934 ( .A(n1259), .Y(n5023) );
  AND2X1 U5935 ( .A(\RF[14][28] ), .B(n10730), .Y(n1247) );
  INVX1 U5936 ( .A(n1247), .Y(n5024) );
  AND2X1 U5937 ( .A(\RF[14][16] ), .B(n10730), .Y(n1235) );
  INVX1 U5938 ( .A(n1235), .Y(n5025) );
  AND2X1 U5939 ( .A(\RF[14][4] ), .B(n10730), .Y(n1223) );
  INVX1 U5940 ( .A(n1223), .Y(n5026) );
  AND2X1 U5941 ( .A(\RF[15][39] ), .B(n10731), .Y(n1192) );
  INVX1 U5942 ( .A(n1192), .Y(n5027) );
  AND2X1 U5943 ( .A(\RF[15][27] ), .B(n10731), .Y(n1180) );
  INVX1 U5944 ( .A(n1180), .Y(n5028) );
  AND2X1 U5945 ( .A(\RF[15][15] ), .B(n10732), .Y(n1168) );
  INVX1 U5946 ( .A(n1168), .Y(n5029) );
  AND2X1 U5947 ( .A(\RF[15][3] ), .B(n10732), .Y(n1156) );
  INVX1 U5948 ( .A(n1156), .Y(n5030) );
  AND2X1 U5949 ( .A(\RF[16][58] ), .B(n10734), .Y(n1146) );
  INVX1 U5950 ( .A(n1146), .Y(n5031) );
  AND2X1 U5951 ( .A(\RF[16][48] ), .B(n10733), .Y(n1136) );
  INVX1 U5952 ( .A(n1136), .Y(n5032) );
  AND2X1 U5953 ( .A(\RF[17][57] ), .B(n10736), .Y(n1080) );
  INVX1 U5954 ( .A(n1080), .Y(n5033) );
  AND2X1 U5955 ( .A(\RF[17][46] ), .B(n10736), .Y(n1069) );
  INVX1 U5956 ( .A(n1069), .Y(n5034) );
  AND2X1 U5957 ( .A(\RF[17][24] ), .B(n10736), .Y(n1047) );
  INVX1 U5958 ( .A(n1047), .Y(n5035) );
  AND2X1 U5959 ( .A(\RF[18][50] ), .B(n10738), .Y(n1008) );
  INVX1 U5960 ( .A(n1008), .Y(n5036) );
  AND2X1 U5961 ( .A(\RF[19][61] ), .B(n10740), .Y(n954) );
  INVX1 U5962 ( .A(n954), .Y(n5037) );
  AND2X1 U5963 ( .A(\RF[19][53] ), .B(n10740), .Y(n946) );
  INVX1 U5964 ( .A(n946), .Y(n5038) );
  AND2X1 U5965 ( .A(\RF[19][49] ), .B(n10740), .Y(n942) );
  INVX1 U5966 ( .A(n942), .Y(n5039) );
  AND2X1 U5967 ( .A(\RF[20][63] ), .B(n10742), .Y(n891) );
  INVX1 U5968 ( .A(n891), .Y(n5040) );
  AND2X1 U5969 ( .A(\RF[20][34] ), .B(n10742), .Y(n862) );
  INVX1 U5970 ( .A(n862), .Y(n5041) );
  AND2X1 U5971 ( .A(\RF[20][22] ), .B(n10741), .Y(n850) );
  INVX1 U5972 ( .A(n850), .Y(n5042) );
  AND2X1 U5973 ( .A(\RF[20][10] ), .B(n10742), .Y(n838) );
  INVX1 U5974 ( .A(n838), .Y(n5043) );
  AND2X1 U5975 ( .A(\RF[21][44] ), .B(n10743), .Y(n807) );
  INVX1 U5976 ( .A(n807), .Y(n5044) );
  AND2X1 U5977 ( .A(\RF[21][33] ), .B(n10744), .Y(n796) );
  INVX1 U5978 ( .A(n796), .Y(n5045) );
  AND2X1 U5979 ( .A(\RF[21][21] ), .B(n10744), .Y(n784) );
  INVX1 U5980 ( .A(n784), .Y(n5046) );
  AND2X1 U5981 ( .A(\RF[21][9] ), .B(n10744), .Y(n772) );
  INVX1 U5982 ( .A(n772), .Y(n5047) );
  AND2X1 U5983 ( .A(\RF[22][59] ), .B(n10746), .Y(n757) );
  INVX1 U5984 ( .A(n757), .Y(n5048) );
  AND2X1 U5985 ( .A(\RF[22][42] ), .B(n10746), .Y(n740) );
  INVX1 U5986 ( .A(n740), .Y(n5049) );
  AND2X1 U5987 ( .A(\RF[22][36] ), .B(n10745), .Y(n734) );
  INVX1 U5988 ( .A(n734), .Y(n5050) );
  AND2X1 U5989 ( .A(\RF[22][12] ), .B(n10745), .Y(n710) );
  INVX1 U5990 ( .A(n710), .Y(n5051) );
  AND2X1 U5991 ( .A(\RF[23][56] ), .B(n10748), .Y(n688) );
  INVX1 U5992 ( .A(n688), .Y(n5052) );
  AND2X1 U5993 ( .A(\RF[23][35] ), .B(n10747), .Y(n667) );
  INVX1 U5994 ( .A(n667), .Y(n5053) );
  AND2X1 U5995 ( .A(\RF[23][23] ), .B(n10748), .Y(n655) );
  INVX1 U5996 ( .A(n655), .Y(n5054) );
  AND2X1 U5997 ( .A(\RF[23][11] ), .B(n10747), .Y(n643) );
  INVX1 U5998 ( .A(n643), .Y(n5055) );
  AND2X1 U5999 ( .A(\RF[24][58] ), .B(n10750), .Y(n623) );
  INVX1 U6000 ( .A(n623), .Y(n5056) );
  AND2X1 U6001 ( .A(\RF[24][48] ), .B(n10749), .Y(n613) );
  INVX1 U6002 ( .A(n613), .Y(n5057) );
  AND2X1 U6003 ( .A(\RF[25][57] ), .B(n10752), .Y(n556) );
  INVX1 U6004 ( .A(n556), .Y(n5058) );
  AND2X1 U6005 ( .A(\RF[25][46] ), .B(n10752), .Y(n545) );
  INVX1 U6006 ( .A(n545), .Y(n5059) );
  AND2X1 U6007 ( .A(\RF[25][24] ), .B(n10752), .Y(n523) );
  INVX1 U6008 ( .A(n523), .Y(n5060) );
  AND2X1 U6009 ( .A(\RF[26][50] ), .B(n10754), .Y(n483) );
  INVX1 U6010 ( .A(n483), .Y(n5061) );
  AND2X1 U6011 ( .A(\RF[27][61] ), .B(n10756), .Y(n428) );
  INVX1 U6012 ( .A(n428), .Y(n5062) );
  AND2X1 U6013 ( .A(\RF[27][53] ), .B(n10756), .Y(n420) );
  INVX1 U6014 ( .A(n420), .Y(n5063) );
  AND2X1 U6015 ( .A(\RF[27][49] ), .B(n10756), .Y(n416) );
  INVX1 U6016 ( .A(n416), .Y(n5064) );
  AND2X1 U6017 ( .A(\RF[28][63] ), .B(n10758), .Y(n364) );
  INVX1 U6018 ( .A(n364), .Y(n5065) );
  AND2X1 U6019 ( .A(\RF[28][34] ), .B(n10758), .Y(n335) );
  INVX1 U6020 ( .A(n335), .Y(n5066) );
  AND2X1 U6021 ( .A(\RF[28][22] ), .B(n10757), .Y(n323) );
  INVX1 U6022 ( .A(n323), .Y(n5067) );
  AND2X1 U6023 ( .A(\RF[28][10] ), .B(n10758), .Y(n311) );
  INVX1 U6024 ( .A(n311), .Y(n5068) );
  AND2X1 U6025 ( .A(\RF[29][44] ), .B(n10759), .Y(n279) );
  INVX1 U6026 ( .A(n279), .Y(n5069) );
  AND2X1 U6027 ( .A(\RF[29][33] ), .B(n10760), .Y(n268) );
  INVX1 U6028 ( .A(n268), .Y(n5070) );
  AND2X1 U6029 ( .A(\RF[29][21] ), .B(n10760), .Y(n256) );
  INVX1 U6030 ( .A(n256), .Y(n5071) );
  AND2X1 U6031 ( .A(\RF[29][9] ), .B(n10760), .Y(n244) );
  INVX1 U6032 ( .A(n244), .Y(n5072) );
  AND2X1 U6033 ( .A(\RF[30][59] ), .B(n10762), .Y(n228) );
  INVX1 U6034 ( .A(n228), .Y(n5073) );
  AND2X1 U6035 ( .A(\RF[30][42] ), .B(n10762), .Y(n211) );
  INVX1 U6036 ( .A(n211), .Y(n5074) );
  AND2X1 U6037 ( .A(\RF[30][36] ), .B(n10761), .Y(n205) );
  INVX1 U6038 ( .A(n205), .Y(n5075) );
  AND2X1 U6039 ( .A(\RF[30][12] ), .B(n10761), .Y(n181) );
  INVX1 U6040 ( .A(n181), .Y(n5076) );
  AND2X1 U6041 ( .A(\RF[31][56] ), .B(n10764), .Y(n151) );
  INVX1 U6042 ( .A(n151), .Y(n5077) );
  AND2X1 U6043 ( .A(\RF[31][35] ), .B(n10763), .Y(n109) );
  INVX1 U6044 ( .A(n109), .Y(n5078) );
  AND2X1 U6045 ( .A(\RF[31][23] ), .B(n10764), .Y(n85) );
  INVX1 U6046 ( .A(n85), .Y(n5079) );
  AND2X1 U6047 ( .A(\RF[31][11] ), .B(n10763), .Y(n61) );
  INVX1 U6048 ( .A(n61), .Y(n5080) );
  AND2X1 U6049 ( .A(\RF[0][39] ), .B(n10702), .Y(n2169) );
  INVX1 U6050 ( .A(n2169), .Y(n5081) );
  AND2X1 U6051 ( .A(\RF[0][27] ), .B(n10702), .Y(n2157) );
  INVX1 U6052 ( .A(n2157), .Y(n5082) );
  AND2X1 U6053 ( .A(\RF[0][15] ), .B(n10701), .Y(n2145) );
  INVX1 U6054 ( .A(n2145), .Y(n5083) );
  AND2X1 U6055 ( .A(\RF[0][3] ), .B(n10702), .Y(n2133) );
  INVX1 U6056 ( .A(n2133), .Y(n5084) );
  AND2X1 U6057 ( .A(\RF[1][40] ), .B(n10704), .Y(n2105) );
  INVX1 U6058 ( .A(n2105), .Y(n5085) );
  AND2X1 U6059 ( .A(\RF[1][28] ), .B(n10704), .Y(n2093) );
  INVX1 U6060 ( .A(n2093), .Y(n5086) );
  AND2X1 U6061 ( .A(\RF[1][16] ), .B(n10703), .Y(n2081) );
  INVX1 U6062 ( .A(n2081), .Y(n5087) );
  AND2X1 U6063 ( .A(\RF[1][4] ), .B(n10704), .Y(n2069) );
  INVX1 U6064 ( .A(n2069), .Y(n5088) );
  AND2X1 U6065 ( .A(\RF[2][45] ), .B(n10706), .Y(n2045) );
  INVX1 U6066 ( .A(n2045), .Y(n5089) );
  AND2X1 U6067 ( .A(\RF[2][32] ), .B(n10706), .Y(n2032) );
  INVX1 U6068 ( .A(n2032), .Y(n5090) );
  AND2X1 U6069 ( .A(\RF[2][13] ), .B(n10705), .Y(n2013) );
  INVX1 U6070 ( .A(n2013), .Y(n5091) );
  AND2X1 U6071 ( .A(\RF[2][1] ), .B(n10706), .Y(n2001) );
  INVX1 U6072 ( .A(n2001), .Y(n5092) );
  AND2X1 U6073 ( .A(\RF[2][0] ), .B(n10706), .Y(n2000) );
  INVX1 U6074 ( .A(n2000), .Y(n5093) );
  AND2X1 U6075 ( .A(\RF[3][37] ), .B(n10708), .Y(n1972) );
  INVX1 U6076 ( .A(n1972), .Y(n5094) );
  AND2X1 U6077 ( .A(\RF[3][26] ), .B(n10708), .Y(n1961) );
  INVX1 U6078 ( .A(n1961), .Y(n5095) );
  AND2X1 U6079 ( .A(\RF[3][14] ), .B(n10708), .Y(n1949) );
  INVX1 U6080 ( .A(n1949), .Y(n5096) );
  AND2X1 U6081 ( .A(\RF[3][2] ), .B(n10708), .Y(n1937) );
  INVX1 U6082 ( .A(n1937), .Y(n5097) );
  AND2X1 U6083 ( .A(\RF[4][61] ), .B(n10710), .Y(n1931) );
  INVX1 U6084 ( .A(n1931), .Y(n5098) );
  AND2X1 U6085 ( .A(\RF[4][53] ), .B(n10710), .Y(n1923) );
  INVX1 U6086 ( .A(n1923), .Y(n5099) );
  AND2X1 U6087 ( .A(\RF[4][49] ), .B(n10710), .Y(n1919) );
  INVX1 U6088 ( .A(n1919), .Y(n5100) );
  AND2X1 U6089 ( .A(\RF[5][50] ), .B(n10712), .Y(n1855) );
  INVX1 U6090 ( .A(n1855), .Y(n5101) );
  AND2X1 U6091 ( .A(\RF[6][57] ), .B(n10714), .Y(n1797) );
  INVX1 U6092 ( .A(n1797), .Y(n5102) );
  AND2X1 U6093 ( .A(\RF[6][46] ), .B(n10714), .Y(n1786) );
  INVX1 U6094 ( .A(n1786), .Y(n5103) );
  AND2X1 U6095 ( .A(\RF[6][24] ), .B(n10714), .Y(n1764) );
  INVX1 U6096 ( .A(n1764), .Y(n5104) );
  AND2X1 U6097 ( .A(\RF[7][58] ), .B(n10716), .Y(n1732) );
  INVX1 U6098 ( .A(n1732), .Y(n5105) );
  AND2X1 U6099 ( .A(\RF[7][48] ), .B(n10716), .Y(n1722) );
  INVX1 U6100 ( .A(n1722), .Y(n5106) );
  AND2X1 U6101 ( .A(\RF[8][56] ), .B(n10718), .Y(n1665) );
  INVX1 U6102 ( .A(n1665), .Y(n5107) );
  AND2X1 U6103 ( .A(\RF[8][35] ), .B(n10717), .Y(n1644) );
  INVX1 U6104 ( .A(n1644), .Y(n5108) );
  AND2X1 U6105 ( .A(\RF[8][23] ), .B(n10718), .Y(n1632) );
  INVX1 U6106 ( .A(n1632), .Y(n5109) );
  AND2X1 U6107 ( .A(\RF[8][11] ), .B(n10718), .Y(n1620) );
  INVX1 U6108 ( .A(n1620), .Y(n5110) );
  AND2X1 U6109 ( .A(\RF[9][59] ), .B(n10720), .Y(n1603) );
  INVX1 U6110 ( .A(n1603), .Y(n5111) );
  AND2X1 U6111 ( .A(\RF[9][42] ), .B(n10720), .Y(n1586) );
  INVX1 U6112 ( .A(n1586), .Y(n5112) );
  AND2X1 U6113 ( .A(\RF[9][36] ), .B(n10719), .Y(n1580) );
  INVX1 U6114 ( .A(n1580), .Y(n5113) );
  AND2X1 U6115 ( .A(\RF[9][12] ), .B(n10720), .Y(n1556) );
  INVX1 U6116 ( .A(n1556), .Y(n5114) );
  AND2X1 U6117 ( .A(\RF[10][44] ), .B(n10722), .Y(n1523) );
  INVX1 U6118 ( .A(n1523), .Y(n5115) );
  AND2X1 U6119 ( .A(\RF[10][33] ), .B(n10722), .Y(n1512) );
  INVX1 U6120 ( .A(n1512), .Y(n5116) );
  AND2X1 U6121 ( .A(\RF[10][21] ), .B(n10722), .Y(n1500) );
  INVX1 U6122 ( .A(n1500), .Y(n5117) );
  AND2X1 U6123 ( .A(\RF[10][9] ), .B(n10722), .Y(n1488) );
  INVX1 U6124 ( .A(n1488), .Y(n5118) );
  AND2X1 U6125 ( .A(\RF[11][63] ), .B(n10724), .Y(n1477) );
  INVX1 U6126 ( .A(n1477), .Y(n5119) );
  AND2X1 U6127 ( .A(\RF[11][34] ), .B(n10724), .Y(n1448) );
  INVX1 U6128 ( .A(n1448), .Y(n5120) );
  AND2X1 U6129 ( .A(\RF[11][22] ), .B(n10724), .Y(n1436) );
  INVX1 U6130 ( .A(n1436), .Y(n5121) );
  AND2X1 U6131 ( .A(\RF[11][10] ), .B(n10724), .Y(n1424) );
  INVX1 U6132 ( .A(n1424), .Y(n5122) );
  AND2X1 U6133 ( .A(\RF[12][39] ), .B(n10726), .Y(n1388) );
  INVX1 U6134 ( .A(n1388), .Y(n5123) );
  AND2X1 U6135 ( .A(\RF[12][27] ), .B(n10726), .Y(n1376) );
  INVX1 U6136 ( .A(n1376), .Y(n5124) );
  AND2X1 U6137 ( .A(\RF[12][15] ), .B(n10725), .Y(n1364) );
  INVX1 U6138 ( .A(n1364), .Y(n5125) );
  AND2X1 U6139 ( .A(\RF[12][3] ), .B(n10726), .Y(n1352) );
  INVX1 U6140 ( .A(n1352), .Y(n5126) );
  AND2X1 U6141 ( .A(\RF[13][40] ), .B(n10728), .Y(n1324) );
  INVX1 U6142 ( .A(n1324), .Y(n5127) );
  AND2X1 U6143 ( .A(\RF[13][28] ), .B(n10728), .Y(n1312) );
  INVX1 U6144 ( .A(n1312), .Y(n5128) );
  AND2X1 U6145 ( .A(\RF[13][16] ), .B(n10727), .Y(n1300) );
  INVX1 U6146 ( .A(n1300), .Y(n5129) );
  AND2X1 U6147 ( .A(\RF[13][4] ), .B(n10728), .Y(n1288) );
  INVX1 U6148 ( .A(n1288), .Y(n5130) );
  AND2X1 U6149 ( .A(\RF[14][45] ), .B(n10730), .Y(n1264) );
  INVX1 U6150 ( .A(n1264), .Y(n5131) );
  AND2X1 U6151 ( .A(\RF[14][32] ), .B(n10730), .Y(n1251) );
  INVX1 U6152 ( .A(n1251), .Y(n5132) );
  AND2X1 U6153 ( .A(\RF[14][13] ), .B(n10729), .Y(n1232) );
  INVX1 U6154 ( .A(n1232), .Y(n5133) );
  AND2X1 U6155 ( .A(\RF[14][1] ), .B(n10730), .Y(n1220) );
  INVX1 U6156 ( .A(n1220), .Y(n5134) );
  AND2X1 U6157 ( .A(\RF[14][0] ), .B(n10730), .Y(n1219) );
  INVX1 U6158 ( .A(n1219), .Y(n5135) );
  AND2X1 U6159 ( .A(\RF[15][37] ), .B(n10732), .Y(n1190) );
  INVX1 U6160 ( .A(n1190), .Y(n5136) );
  AND2X1 U6161 ( .A(\RF[15][26] ), .B(n10732), .Y(n1179) );
  INVX1 U6162 ( .A(n1179), .Y(n5137) );
  AND2X1 U6163 ( .A(\RF[15][14] ), .B(n10732), .Y(n1167) );
  INVX1 U6164 ( .A(n1167), .Y(n5138) );
  AND2X1 U6165 ( .A(\RF[15][2] ), .B(n10732), .Y(n1155) );
  INVX1 U6166 ( .A(n1155), .Y(n5139) );
  AND2X1 U6167 ( .A(\RF[16][61] ), .B(n10734), .Y(n1149) );
  INVX1 U6168 ( .A(n1149), .Y(n5140) );
  AND2X1 U6169 ( .A(\RF[16][53] ), .B(n10734), .Y(n1141) );
  INVX1 U6170 ( .A(n1141), .Y(n5141) );
  AND2X1 U6171 ( .A(\RF[16][49] ), .B(n10734), .Y(n1137) );
  INVX1 U6172 ( .A(n1137), .Y(n5142) );
  AND2X1 U6173 ( .A(\RF[17][50] ), .B(n10736), .Y(n1073) );
  INVX1 U6174 ( .A(n1073), .Y(n5143) );
  AND2X1 U6175 ( .A(\RF[18][57] ), .B(n10738), .Y(n1015) );
  INVX1 U6176 ( .A(n1015), .Y(n5144) );
  AND2X1 U6177 ( .A(\RF[18][46] ), .B(n10738), .Y(n1004) );
  INVX1 U6178 ( .A(n1004), .Y(n5145) );
  AND2X1 U6179 ( .A(\RF[18][24] ), .B(n10738), .Y(n982) );
  INVX1 U6180 ( .A(n982), .Y(n5146) );
  AND2X1 U6181 ( .A(\RF[19][58] ), .B(n10740), .Y(n951) );
  INVX1 U6182 ( .A(n951), .Y(n5147) );
  AND2X1 U6183 ( .A(\RF[19][48] ), .B(n10740), .Y(n941) );
  INVX1 U6184 ( .A(n941), .Y(n5148) );
  AND2X1 U6185 ( .A(\RF[20][56] ), .B(n10742), .Y(n884) );
  INVX1 U6186 ( .A(n884), .Y(n5149) );
  AND2X1 U6187 ( .A(\RF[20][35] ), .B(n10741), .Y(n863) );
  INVX1 U6188 ( .A(n863), .Y(n5150) );
  AND2X1 U6189 ( .A(\RF[20][23] ), .B(n10742), .Y(n851) );
  INVX1 U6190 ( .A(n851), .Y(n5151) );
  AND2X1 U6191 ( .A(\RF[20][11] ), .B(n10742), .Y(n839) );
  INVX1 U6192 ( .A(n839), .Y(n5152) );
  AND2X1 U6193 ( .A(\RF[21][59] ), .B(n10744), .Y(n822) );
  INVX1 U6194 ( .A(n822), .Y(n5153) );
  AND2X1 U6195 ( .A(\RF[21][42] ), .B(n10744), .Y(n805) );
  INVX1 U6196 ( .A(n805), .Y(n5154) );
  AND2X1 U6197 ( .A(\RF[21][36] ), .B(n10743), .Y(n799) );
  INVX1 U6198 ( .A(n799), .Y(n5155) );
  AND2X1 U6199 ( .A(\RF[21][12] ), .B(n10744), .Y(n775) );
  INVX1 U6200 ( .A(n775), .Y(n5156) );
  AND2X1 U6201 ( .A(\RF[22][44] ), .B(n10746), .Y(n742) );
  INVX1 U6202 ( .A(n742), .Y(n5157) );
  AND2X1 U6203 ( .A(\RF[22][33] ), .B(n10746), .Y(n731) );
  INVX1 U6204 ( .A(n731), .Y(n5158) );
  AND2X1 U6205 ( .A(\RF[22][21] ), .B(n10746), .Y(n719) );
  INVX1 U6206 ( .A(n719), .Y(n5159) );
  AND2X1 U6207 ( .A(\RF[22][9] ), .B(n10746), .Y(n707) );
  INVX1 U6208 ( .A(n707), .Y(n5160) );
  AND2X1 U6209 ( .A(\RF[23][63] ), .B(n10748), .Y(n695) );
  INVX1 U6210 ( .A(n695), .Y(n5161) );
  AND2X1 U6211 ( .A(\RF[23][34] ), .B(n10748), .Y(n666) );
  INVX1 U6212 ( .A(n666), .Y(n5162) );
  AND2X1 U6213 ( .A(\RF[23][22] ), .B(n10748), .Y(n654) );
  INVX1 U6214 ( .A(n654), .Y(n5163) );
  AND2X1 U6215 ( .A(\RF[23][10] ), .B(n10748), .Y(n642) );
  INVX1 U6216 ( .A(n642), .Y(n5164) );
  AND2X1 U6217 ( .A(\RF[24][61] ), .B(n10750), .Y(n626) );
  INVX1 U6218 ( .A(n626), .Y(n5165) );
  AND2X1 U6219 ( .A(\RF[24][53] ), .B(n10750), .Y(n618) );
  INVX1 U6220 ( .A(n618), .Y(n5166) );
  AND2X1 U6221 ( .A(\RF[24][49] ), .B(n10750), .Y(n614) );
  INVX1 U6222 ( .A(n614), .Y(n5167) );
  AND2X1 U6223 ( .A(\RF[25][50] ), .B(n10752), .Y(n549) );
  INVX1 U6224 ( .A(n549), .Y(n5168) );
  AND2X1 U6225 ( .A(\RF[26][57] ), .B(n10754), .Y(n490) );
  INVX1 U6226 ( .A(n490), .Y(n5169) );
  AND2X1 U6227 ( .A(\RF[26][46] ), .B(n10754), .Y(n479) );
  INVX1 U6228 ( .A(n479), .Y(n5170) );
  AND2X1 U6229 ( .A(\RF[26][24] ), .B(n10754), .Y(n457) );
  INVX1 U6230 ( .A(n457), .Y(n5171) );
  AND2X1 U6231 ( .A(\RF[27][58] ), .B(n10756), .Y(n425) );
  INVX1 U6232 ( .A(n425), .Y(n5172) );
  AND2X1 U6233 ( .A(\RF[27][48] ), .B(n10756), .Y(n415) );
  INVX1 U6234 ( .A(n415), .Y(n5173) );
  AND2X1 U6235 ( .A(\RF[28][56] ), .B(n10758), .Y(n357) );
  INVX1 U6236 ( .A(n357), .Y(n5174) );
  AND2X1 U6237 ( .A(\RF[28][35] ), .B(n10757), .Y(n336) );
  INVX1 U6238 ( .A(n336), .Y(n5175) );
  AND2X1 U6239 ( .A(\RF[28][23] ), .B(n10758), .Y(n324) );
  INVX1 U6240 ( .A(n324), .Y(n5176) );
  AND2X1 U6241 ( .A(\RF[28][11] ), .B(n10758), .Y(n312) );
  INVX1 U6242 ( .A(n312), .Y(n5177) );
  AND2X1 U6243 ( .A(\RF[29][59] ), .B(n10760), .Y(n294) );
  INVX1 U6244 ( .A(n294), .Y(n5178) );
  AND2X1 U6245 ( .A(\RF[29][42] ), .B(n10760), .Y(n277) );
  INVX1 U6246 ( .A(n277), .Y(n5179) );
  AND2X1 U6247 ( .A(\RF[29][36] ), .B(n10759), .Y(n271) );
  INVX1 U6248 ( .A(n271), .Y(n5180) );
  AND2X1 U6249 ( .A(\RF[29][12] ), .B(n10760), .Y(n247) );
  INVX1 U6250 ( .A(n247), .Y(n5181) );
  AND2X1 U6251 ( .A(\RF[30][44] ), .B(n10762), .Y(n213) );
  INVX1 U6252 ( .A(n213), .Y(n5182) );
  AND2X1 U6253 ( .A(\RF[30][33] ), .B(n10762), .Y(n202) );
  INVX1 U6254 ( .A(n202), .Y(n5183) );
  AND2X1 U6255 ( .A(\RF[30][21] ), .B(n10762), .Y(n190) );
  INVX1 U6256 ( .A(n190), .Y(n5184) );
  AND2X1 U6257 ( .A(\RF[30][9] ), .B(n10762), .Y(n178) );
  INVX1 U6258 ( .A(n178), .Y(n5185) );
  AND2X1 U6259 ( .A(\RF[31][63] ), .B(n10764), .Y(n165) );
  INVX1 U6260 ( .A(n165), .Y(n5186) );
  AND2X1 U6261 ( .A(\RF[31][34] ), .B(n10764), .Y(n107) );
  INVX1 U6262 ( .A(n107), .Y(n5187) );
  AND2X1 U6263 ( .A(\RF[31][22] ), .B(n10764), .Y(n83) );
  INVX1 U6264 ( .A(n83), .Y(n5188) );
  AND2X1 U6265 ( .A(\RF[31][10] ), .B(n10764), .Y(n59) );
  INVX1 U6266 ( .A(n59), .Y(n5189) );
  AND2X1 U6267 ( .A(\RF[0][40] ), .B(n10701), .Y(n2170) );
  INVX1 U6268 ( .A(n2170), .Y(n5190) );
  AND2X1 U6269 ( .A(\RF[0][28] ), .B(n10702), .Y(n2158) );
  INVX1 U6270 ( .A(n2158), .Y(n5191) );
  AND2X1 U6271 ( .A(\RF[0][16] ), .B(n10702), .Y(n2146) );
  INVX1 U6272 ( .A(n2146), .Y(n5192) );
  AND2X1 U6273 ( .A(\RF[0][4] ), .B(n10702), .Y(n2134) );
  INVX1 U6274 ( .A(n2134), .Y(n5193) );
  AND2X1 U6275 ( .A(\RF[1][39] ), .B(n10703), .Y(n2104) );
  INVX1 U6276 ( .A(n2104), .Y(n5194) );
  AND2X1 U6277 ( .A(\RF[1][27] ), .B(n10704), .Y(n2092) );
  INVX1 U6278 ( .A(n2092), .Y(n5195) );
  AND2X1 U6279 ( .A(\RF[1][15] ), .B(n10704), .Y(n2080) );
  INVX1 U6280 ( .A(n2080), .Y(n5196) );
  AND2X1 U6281 ( .A(\RF[1][3] ), .B(n10704), .Y(n2068) );
  INVX1 U6282 ( .A(n2068), .Y(n5197) );
  AND2X1 U6283 ( .A(\RF[2][37] ), .B(n10705), .Y(n2037) );
  INVX1 U6284 ( .A(n2037), .Y(n5198) );
  AND2X1 U6285 ( .A(\RF[2][26] ), .B(n10706), .Y(n2026) );
  INVX1 U6286 ( .A(n2026), .Y(n5199) );
  AND2X1 U6287 ( .A(\RF[2][14] ), .B(n10706), .Y(n2014) );
  INVX1 U6288 ( .A(n2014), .Y(n5200) );
  AND2X1 U6289 ( .A(\RF[2][2] ), .B(n10706), .Y(n2002) );
  INVX1 U6290 ( .A(n2002), .Y(n5201) );
  AND2X1 U6291 ( .A(\RF[3][45] ), .B(n10708), .Y(n1980) );
  INVX1 U6292 ( .A(n1980), .Y(n5202) );
  AND2X1 U6293 ( .A(\RF[3][32] ), .B(n10707), .Y(n1967) );
  INVX1 U6294 ( .A(n1967), .Y(n5203) );
  AND2X1 U6295 ( .A(\RF[3][13] ), .B(n10708), .Y(n1948) );
  INVX1 U6296 ( .A(n1948), .Y(n5204) );
  AND2X1 U6297 ( .A(\RF[3][1] ), .B(n10707), .Y(n1936) );
  INVX1 U6298 ( .A(n1936), .Y(n5205) );
  AND2X1 U6299 ( .A(\RF[3][0] ), .B(n10708), .Y(n1935) );
  INVX1 U6300 ( .A(n1935), .Y(n5206) );
  AND2X1 U6301 ( .A(\RF[4][50] ), .B(n10710), .Y(n1920) );
  INVX1 U6302 ( .A(n1920), .Y(n5207) );
  AND2X1 U6303 ( .A(\RF[5][61] ), .B(n10712), .Y(n1866) );
  INVX1 U6304 ( .A(n1866), .Y(n5208) );
  AND2X1 U6305 ( .A(\RF[5][53] ), .B(n10712), .Y(n1858) );
  INVX1 U6306 ( .A(n1858), .Y(n5209) );
  AND2X1 U6307 ( .A(\RF[5][49] ), .B(n10712), .Y(n1854) );
  INVX1 U6308 ( .A(n1854), .Y(n5210) );
  AND2X1 U6309 ( .A(\RF[6][58] ), .B(n10714), .Y(n1798) );
  INVX1 U6310 ( .A(n1798), .Y(n5211) );
  AND2X1 U6311 ( .A(\RF[6][48] ), .B(n10714), .Y(n1788) );
  INVX1 U6312 ( .A(n1788), .Y(n5212) );
  AND2X1 U6313 ( .A(\RF[7][57] ), .B(n10716), .Y(n1731) );
  INVX1 U6314 ( .A(n1731), .Y(n5213) );
  AND2X1 U6315 ( .A(\RF[7][46] ), .B(n10716), .Y(n1720) );
  INVX1 U6316 ( .A(n1720), .Y(n5214) );
  AND2X1 U6317 ( .A(\RF[7][24] ), .B(n10716), .Y(n1698) );
  INVX1 U6318 ( .A(n1698), .Y(n5215) );
  AND2X1 U6319 ( .A(\RF[8][59] ), .B(n10718), .Y(n1668) );
  INVX1 U6320 ( .A(n1668), .Y(n5216) );
  AND2X1 U6321 ( .A(\RF[8][42] ), .B(n10718), .Y(n1651) );
  INVX1 U6322 ( .A(n1651), .Y(n5217) );
  AND2X1 U6323 ( .A(\RF[8][36] ), .B(n10718), .Y(n1645) );
  INVX1 U6324 ( .A(n1645), .Y(n5218) );
  AND2X1 U6325 ( .A(\RF[8][12] ), .B(n10718), .Y(n1621) );
  INVX1 U6326 ( .A(n1621), .Y(n5219) );
  AND2X1 U6327 ( .A(\RF[9][56] ), .B(n10720), .Y(n1600) );
  INVX1 U6328 ( .A(n1600), .Y(n5220) );
  AND2X1 U6329 ( .A(\RF[9][35] ), .B(n10720), .Y(n1579) );
  INVX1 U6330 ( .A(n1579), .Y(n5221) );
  AND2X1 U6331 ( .A(\RF[9][23] ), .B(n10720), .Y(n1567) );
  INVX1 U6332 ( .A(n1567), .Y(n5222) );
  AND2X1 U6333 ( .A(\RF[9][11] ), .B(n10720), .Y(n1555) );
  INVX1 U6334 ( .A(n1555), .Y(n5223) );
  AND2X1 U6335 ( .A(\RF[10][63] ), .B(n10722), .Y(n1542) );
  INVX1 U6336 ( .A(n1542), .Y(n5224) );
  AND2X1 U6337 ( .A(\RF[10][34] ), .B(n10722), .Y(n1513) );
  INVX1 U6338 ( .A(n1513), .Y(n5225) );
  AND2X1 U6339 ( .A(\RF[10][22] ), .B(n10722), .Y(n1501) );
  INVX1 U6340 ( .A(n1501), .Y(n5226) );
  AND2X1 U6341 ( .A(\RF[10][10] ), .B(n10722), .Y(n1489) );
  INVX1 U6342 ( .A(n1489), .Y(n5227) );
  AND2X1 U6343 ( .A(\RF[11][44] ), .B(n10724), .Y(n1458) );
  INVX1 U6344 ( .A(n1458), .Y(n5228) );
  AND2X1 U6345 ( .A(\RF[11][33] ), .B(n10724), .Y(n1447) );
  INVX1 U6346 ( .A(n1447), .Y(n5229) );
  AND2X1 U6347 ( .A(\RF[11][21] ), .B(n10724), .Y(n1435) );
  INVX1 U6348 ( .A(n1435), .Y(n5230) );
  AND2X1 U6349 ( .A(\RF[11][9] ), .B(n10724), .Y(n1423) );
  INVX1 U6350 ( .A(n1423), .Y(n5231) );
  AND2X1 U6351 ( .A(\RF[12][40] ), .B(n10725), .Y(n1389) );
  INVX1 U6352 ( .A(n1389), .Y(n5232) );
  AND2X1 U6353 ( .A(\RF[12][28] ), .B(n10726), .Y(n1377) );
  INVX1 U6354 ( .A(n1377), .Y(n5233) );
  AND2X1 U6355 ( .A(\RF[12][16] ), .B(n10726), .Y(n1365) );
  INVX1 U6356 ( .A(n1365), .Y(n5234) );
  AND2X1 U6357 ( .A(\RF[12][4] ), .B(n10726), .Y(n1353) );
  INVX1 U6358 ( .A(n1353), .Y(n5235) );
  AND2X1 U6359 ( .A(\RF[13][39] ), .B(n10727), .Y(n1323) );
  INVX1 U6360 ( .A(n1323), .Y(n5236) );
  AND2X1 U6361 ( .A(\RF[13][27] ), .B(n10728), .Y(n1311) );
  INVX1 U6362 ( .A(n1311), .Y(n5237) );
  AND2X1 U6363 ( .A(\RF[13][15] ), .B(n10728), .Y(n1299) );
  INVX1 U6364 ( .A(n1299), .Y(n5238) );
  AND2X1 U6365 ( .A(\RF[13][3] ), .B(n10728), .Y(n1287) );
  INVX1 U6366 ( .A(n1287), .Y(n5239) );
  AND2X1 U6367 ( .A(\RF[14][37] ), .B(n10729), .Y(n1256) );
  INVX1 U6368 ( .A(n1256), .Y(n5240) );
  AND2X1 U6369 ( .A(\RF[14][26] ), .B(n10730), .Y(n1245) );
  INVX1 U6370 ( .A(n1245), .Y(n5241) );
  AND2X1 U6371 ( .A(\RF[14][14] ), .B(n10730), .Y(n1233) );
  INVX1 U6372 ( .A(n1233), .Y(n5242) );
  AND2X1 U6373 ( .A(\RF[14][2] ), .B(n10730), .Y(n1221) );
  INVX1 U6374 ( .A(n1221), .Y(n5243) );
  AND2X1 U6375 ( .A(\RF[15][45] ), .B(n10732), .Y(n1198) );
  INVX1 U6376 ( .A(n1198), .Y(n5244) );
  AND2X1 U6377 ( .A(\RF[15][32] ), .B(n10731), .Y(n1185) );
  INVX1 U6378 ( .A(n1185), .Y(n5245) );
  AND2X1 U6379 ( .A(\RF[15][13] ), .B(n10732), .Y(n1166) );
  INVX1 U6380 ( .A(n1166), .Y(n5246) );
  AND2X1 U6381 ( .A(\RF[15][1] ), .B(n10731), .Y(n1154) );
  INVX1 U6382 ( .A(n1154), .Y(n5247) );
  AND2X1 U6383 ( .A(\RF[15][0] ), .B(n10732), .Y(n1153) );
  INVX1 U6384 ( .A(n1153), .Y(n5248) );
  AND2X1 U6385 ( .A(\RF[16][50] ), .B(n10734), .Y(n1138) );
  INVX1 U6386 ( .A(n1138), .Y(n5249) );
  AND2X1 U6387 ( .A(\RF[17][61] ), .B(n10736), .Y(n1084) );
  INVX1 U6388 ( .A(n1084), .Y(n5250) );
  AND2X1 U6389 ( .A(\RF[17][53] ), .B(n10736), .Y(n1076) );
  INVX1 U6390 ( .A(n1076), .Y(n5251) );
  AND2X1 U6391 ( .A(\RF[17][49] ), .B(n10736), .Y(n1072) );
  INVX1 U6392 ( .A(n1072), .Y(n5252) );
  AND2X1 U6393 ( .A(\RF[18][58] ), .B(n10738), .Y(n1016) );
  INVX1 U6394 ( .A(n1016), .Y(n5253) );
  AND2X1 U6395 ( .A(\RF[18][48] ), .B(n10738), .Y(n1006) );
  INVX1 U6396 ( .A(n1006), .Y(n5254) );
  AND2X1 U6397 ( .A(\RF[19][57] ), .B(n10740), .Y(n950) );
  INVX1 U6398 ( .A(n950), .Y(n5255) );
  AND2X1 U6399 ( .A(\RF[19][46] ), .B(n10740), .Y(n939) );
  INVX1 U6400 ( .A(n939), .Y(n5256) );
  AND2X1 U6401 ( .A(\RF[19][24] ), .B(n10740), .Y(n917) );
  INVX1 U6402 ( .A(n917), .Y(n5257) );
  AND2X1 U6403 ( .A(\RF[20][59] ), .B(n10742), .Y(n887) );
  INVX1 U6404 ( .A(n887), .Y(n5258) );
  AND2X1 U6405 ( .A(\RF[20][42] ), .B(n10742), .Y(n870) );
  INVX1 U6406 ( .A(n870), .Y(n5259) );
  AND2X1 U6407 ( .A(\RF[20][36] ), .B(n10742), .Y(n864) );
  INVX1 U6408 ( .A(n864), .Y(n5260) );
  AND2X1 U6409 ( .A(\RF[20][12] ), .B(n10742), .Y(n840) );
  INVX1 U6410 ( .A(n840), .Y(n5261) );
  AND2X1 U6411 ( .A(\RF[21][56] ), .B(n10744), .Y(n819) );
  INVX1 U6412 ( .A(n819), .Y(n5262) );
  AND2X1 U6413 ( .A(\RF[21][35] ), .B(n10744), .Y(n798) );
  INVX1 U6414 ( .A(n798), .Y(n5263) );
  AND2X1 U6415 ( .A(\RF[21][23] ), .B(n10744), .Y(n786) );
  INVX1 U6416 ( .A(n786), .Y(n5264) );
  AND2X1 U6417 ( .A(\RF[21][11] ), .B(n10744), .Y(n774) );
  INVX1 U6418 ( .A(n774), .Y(n5265) );
  AND2X1 U6419 ( .A(\RF[22][63] ), .B(n10746), .Y(n761) );
  INVX1 U6420 ( .A(n761), .Y(n5266) );
  AND2X1 U6421 ( .A(\RF[22][34] ), .B(n10746), .Y(n732) );
  INVX1 U6422 ( .A(n732), .Y(n5267) );
  AND2X1 U6423 ( .A(\RF[22][22] ), .B(n10746), .Y(n720) );
  INVX1 U6424 ( .A(n720), .Y(n5268) );
  AND2X1 U6425 ( .A(\RF[22][10] ), .B(n10746), .Y(n708) );
  INVX1 U6426 ( .A(n708), .Y(n5269) );
  AND2X1 U6427 ( .A(\RF[23][44] ), .B(n10748), .Y(n676) );
  INVX1 U6428 ( .A(n676), .Y(n5270) );
  AND2X1 U6429 ( .A(\RF[23][33] ), .B(n10748), .Y(n665) );
  INVX1 U6430 ( .A(n665), .Y(n5271) );
  AND2X1 U6431 ( .A(\RF[23][21] ), .B(n10748), .Y(n653) );
  INVX1 U6432 ( .A(n653), .Y(n5272) );
  AND2X1 U6433 ( .A(\RF[23][9] ), .B(n10748), .Y(n641) );
  INVX1 U6434 ( .A(n641), .Y(n5273) );
  AND2X1 U6435 ( .A(\RF[24][50] ), .B(n10750), .Y(n615) );
  INVX1 U6436 ( .A(n615), .Y(n5274) );
  AND2X1 U6437 ( .A(\RF[25][61] ), .B(n10752), .Y(n560) );
  INVX1 U6438 ( .A(n560), .Y(n5275) );
  AND2X1 U6439 ( .A(\RF[25][53] ), .B(n10752), .Y(n552) );
  INVX1 U6440 ( .A(n552), .Y(n5276) );
  AND2X1 U6441 ( .A(\RF[25][49] ), .B(n10752), .Y(n548) );
  INVX1 U6442 ( .A(n548), .Y(n5277) );
  AND2X1 U6443 ( .A(\RF[26][58] ), .B(n10754), .Y(n491) );
  INVX1 U6444 ( .A(n491), .Y(n5278) );
  AND2X1 U6445 ( .A(\RF[26][48] ), .B(n10754), .Y(n481) );
  INVX1 U6446 ( .A(n481), .Y(n5279) );
  AND2X1 U6447 ( .A(\RF[27][57] ), .B(n10756), .Y(n424) );
  INVX1 U6448 ( .A(n424), .Y(n5280) );
  AND2X1 U6449 ( .A(\RF[27][46] ), .B(n10756), .Y(n413) );
  INVX1 U6450 ( .A(n413), .Y(n5281) );
  AND2X1 U6451 ( .A(\RF[27][24] ), .B(n10756), .Y(n391) );
  INVX1 U6452 ( .A(n391), .Y(n5282) );
  AND2X1 U6453 ( .A(\RF[28][59] ), .B(n10758), .Y(n360) );
  INVX1 U6454 ( .A(n360), .Y(n5283) );
  AND2X1 U6455 ( .A(\RF[28][42] ), .B(n10758), .Y(n343) );
  INVX1 U6456 ( .A(n343), .Y(n5284) );
  AND2X1 U6457 ( .A(\RF[28][36] ), .B(n10758), .Y(n337) );
  INVX1 U6458 ( .A(n337), .Y(n5285) );
  AND2X1 U6459 ( .A(\RF[28][12] ), .B(n10758), .Y(n313) );
  INVX1 U6460 ( .A(n313), .Y(n5286) );
  AND2X1 U6461 ( .A(\RF[29][56] ), .B(n10760), .Y(n291) );
  INVX1 U6462 ( .A(n291), .Y(n5287) );
  AND2X1 U6463 ( .A(\RF[29][35] ), .B(n10760), .Y(n270) );
  INVX1 U6464 ( .A(n270), .Y(n5288) );
  AND2X1 U6465 ( .A(\RF[29][23] ), .B(n10760), .Y(n258) );
  INVX1 U6466 ( .A(n258), .Y(n5289) );
  AND2X1 U6467 ( .A(\RF[29][11] ), .B(n10760), .Y(n246) );
  INVX1 U6468 ( .A(n246), .Y(n5290) );
  AND2X1 U6469 ( .A(\RF[30][63] ), .B(n10762), .Y(n232) );
  INVX1 U6470 ( .A(n232), .Y(n5291) );
  AND2X1 U6471 ( .A(\RF[30][34] ), .B(n10762), .Y(n203) );
  INVX1 U6472 ( .A(n203), .Y(n5292) );
  AND2X1 U6473 ( .A(\RF[30][22] ), .B(n10762), .Y(n191) );
  INVX1 U6474 ( .A(n191), .Y(n5293) );
  AND2X1 U6475 ( .A(\RF[30][10] ), .B(n10762), .Y(n179) );
  INVX1 U6476 ( .A(n179), .Y(n5294) );
  AND2X1 U6477 ( .A(\RF[31][44] ), .B(n10764), .Y(n127) );
  INVX1 U6478 ( .A(n127), .Y(n5295) );
  AND2X1 U6479 ( .A(\RF[31][33] ), .B(n10764), .Y(n105) );
  INVX1 U6480 ( .A(n105), .Y(n5296) );
  AND2X1 U6481 ( .A(\RF[31][21] ), .B(n10764), .Y(n81) );
  INVX1 U6482 ( .A(n81), .Y(n5297) );
  AND2X1 U6483 ( .A(\RF[31][9] ), .B(n10764), .Y(n57) );
  INVX1 U6484 ( .A(n57), .Y(n5298) );
  BUFX2 U6485 ( .A(n630), .Y(n5299) );
  AND2X1 U6486 ( .A(\RF[0][57] ), .B(n10702), .Y(n2187) );
  INVX1 U6487 ( .A(n2187), .Y(n5300) );
  AND2X1 U6488 ( .A(\RF[0][46] ), .B(n10701), .Y(n2176) );
  INVX1 U6489 ( .A(n2176), .Y(n5301) );
  AND2X1 U6490 ( .A(\RF[0][24] ), .B(n10701), .Y(n2154) );
  INVX1 U6491 ( .A(n2154), .Y(n5302) );
  AND2X1 U6492 ( .A(\RF[1][58] ), .B(n10704), .Y(n2123) );
  INVX1 U6493 ( .A(n2123), .Y(n5303) );
  AND2X1 U6494 ( .A(\RF[1][48] ), .B(n10703), .Y(n2113) );
  INVX1 U6495 ( .A(n2113), .Y(n5304) );
  AND2X1 U6496 ( .A(\RF[2][61] ), .B(n10706), .Y(n2061) );
  INVX1 U6497 ( .A(n2061), .Y(n5305) );
  AND2X1 U6498 ( .A(\RF[2][53] ), .B(n10706), .Y(n2053) );
  INVX1 U6499 ( .A(n2053), .Y(n5306) );
  AND2X1 U6500 ( .A(\RF[2][49] ), .B(n10705), .Y(n2049) );
  INVX1 U6501 ( .A(n2049), .Y(n5307) );
  AND2X1 U6502 ( .A(\RF[3][50] ), .B(n10707), .Y(n1985) );
  INVX1 U6503 ( .A(n1985), .Y(n5308) );
  AND2X1 U6504 ( .A(\RF[4][45] ), .B(n10709), .Y(n1915) );
  INVX1 U6505 ( .A(n1915), .Y(n5309) );
  AND2X1 U6506 ( .A(\RF[4][32] ), .B(n10709), .Y(n1902) );
  INVX1 U6507 ( .A(n1902), .Y(n5310) );
  AND2X1 U6508 ( .A(\RF[4][13] ), .B(n10710), .Y(n1883) );
  INVX1 U6509 ( .A(n1883), .Y(n5311) );
  AND2X1 U6510 ( .A(\RF[4][1] ), .B(n10709), .Y(n1871) );
  INVX1 U6511 ( .A(n1871), .Y(n5312) );
  AND2X1 U6512 ( .A(\RF[4][0] ), .B(n10709), .Y(n1870) );
  INVX1 U6513 ( .A(n1870), .Y(n5313) );
  AND2X1 U6514 ( .A(\RF[5][37] ), .B(n10711), .Y(n1842) );
  INVX1 U6515 ( .A(n1842), .Y(n5314) );
  AND2X1 U6516 ( .A(\RF[5][26] ), .B(n10712), .Y(n1831) );
  INVX1 U6517 ( .A(n1831), .Y(n5315) );
  AND2X1 U6518 ( .A(\RF[5][14] ), .B(n10711), .Y(n1819) );
  INVX1 U6519 ( .A(n1819), .Y(n5316) );
  AND2X1 U6520 ( .A(\RF[5][2] ), .B(n10712), .Y(n1807) );
  INVX1 U6521 ( .A(n1807), .Y(n5317) );
  AND2X1 U6522 ( .A(\RF[6][39] ), .B(n10713), .Y(n1779) );
  INVX1 U6523 ( .A(n1779), .Y(n5318) );
  AND2X1 U6524 ( .A(\RF[6][27] ), .B(n10714), .Y(n1767) );
  INVX1 U6525 ( .A(n1767), .Y(n5319) );
  AND2X1 U6526 ( .A(\RF[6][15] ), .B(n10713), .Y(n1755) );
  INVX1 U6527 ( .A(n1755), .Y(n5320) );
  AND2X1 U6528 ( .A(\RF[6][3] ), .B(n10714), .Y(n1743) );
  INVX1 U6529 ( .A(n1743), .Y(n5321) );
  AND2X1 U6530 ( .A(\RF[7][40] ), .B(n10715), .Y(n1714) );
  INVX1 U6531 ( .A(n1714), .Y(n5322) );
  AND2X1 U6532 ( .A(\RF[7][28] ), .B(n10716), .Y(n1702) );
  INVX1 U6533 ( .A(n1702), .Y(n5323) );
  AND2X1 U6534 ( .A(\RF[7][16] ), .B(n10715), .Y(n1690) );
  INVX1 U6535 ( .A(n1690), .Y(n5324) );
  AND2X1 U6536 ( .A(\RF[7][4] ), .B(n10716), .Y(n1678) );
  INVX1 U6537 ( .A(n1678), .Y(n5325) );
  AND2X1 U6538 ( .A(\RF[8][41] ), .B(n10717), .Y(n1650) );
  INVX1 U6539 ( .A(n1650), .Y(n5326) );
  AND2X1 U6540 ( .A(\RF[8][29] ), .B(n10718), .Y(n1638) );
  INVX1 U6541 ( .A(n1638), .Y(n5327) );
  AND2X1 U6542 ( .A(\RF[8][17] ), .B(n10717), .Y(n1626) );
  INVX1 U6543 ( .A(n1626), .Y(n5328) );
  AND2X1 U6544 ( .A(\RF[8][5] ), .B(n10718), .Y(n1614) );
  INVX1 U6545 ( .A(n1614), .Y(n5329) );
  AND2X1 U6546 ( .A(\RF[9][38] ), .B(n10720), .Y(n1582) );
  INVX1 U6547 ( .A(n1582), .Y(n5330) );
  AND2X1 U6548 ( .A(\RF[9][30] ), .B(n10719), .Y(n1574) );
  INVX1 U6549 ( .A(n1574), .Y(n5331) );
  AND2X1 U6550 ( .A(\RF[9][18] ), .B(n10719), .Y(n1562) );
  INVX1 U6551 ( .A(n1562), .Y(n5332) );
  AND2X1 U6552 ( .A(\RF[9][6] ), .B(n10720), .Y(n1550) );
  INVX1 U6553 ( .A(n1550), .Y(n5333) );
  AND2X1 U6554 ( .A(\RF[10][43] ), .B(n10721), .Y(n1522) );
  INVX1 U6555 ( .A(n1522), .Y(n5334) );
  AND2X1 U6556 ( .A(\RF[10][31] ), .B(n10722), .Y(n1510) );
  INVX1 U6557 ( .A(n1510), .Y(n5335) );
  AND2X1 U6558 ( .A(\RF[10][19] ), .B(n10721), .Y(n1498) );
  INVX1 U6559 ( .A(n1498), .Y(n5336) );
  AND2X1 U6560 ( .A(\RF[10][7] ), .B(n10722), .Y(n1486) );
  INVX1 U6561 ( .A(n1486), .Y(n5337) );
  AND2X1 U6562 ( .A(\RF[11][47] ), .B(n10723), .Y(n1461) );
  INVX1 U6563 ( .A(n1461), .Y(n5338) );
  AND2X1 U6564 ( .A(\RF[11][25] ), .B(n10723), .Y(n1439) );
  INVX1 U6565 ( .A(n1439), .Y(n5339) );
  AND2X1 U6566 ( .A(\RF[11][20] ), .B(n10724), .Y(n1434) );
  INVX1 U6567 ( .A(n1434), .Y(n5340) );
  AND2X1 U6568 ( .A(\RF[11][8] ), .B(n10724), .Y(n1422) );
  INVX1 U6569 ( .A(n1422), .Y(n5341) );
  AND2X1 U6570 ( .A(\RF[12][57] ), .B(n10726), .Y(n1406) );
  INVX1 U6571 ( .A(n1406), .Y(n5342) );
  AND2X1 U6572 ( .A(\RF[12][46] ), .B(n10725), .Y(n1395) );
  INVX1 U6573 ( .A(n1395), .Y(n5343) );
  AND2X1 U6574 ( .A(\RF[12][24] ), .B(n10725), .Y(n1373) );
  INVX1 U6575 ( .A(n1373), .Y(n5344) );
  AND2X1 U6576 ( .A(\RF[13][58] ), .B(n10728), .Y(n1342) );
  INVX1 U6577 ( .A(n1342), .Y(n5345) );
  AND2X1 U6578 ( .A(\RF[13][48] ), .B(n10727), .Y(n1332) );
  INVX1 U6579 ( .A(n1332), .Y(n5346) );
  AND2X1 U6580 ( .A(\RF[14][61] ), .B(n10730), .Y(n1280) );
  INVX1 U6581 ( .A(n1280), .Y(n5347) );
  AND2X1 U6582 ( .A(\RF[14][53] ), .B(n10730), .Y(n1272) );
  INVX1 U6583 ( .A(n1272), .Y(n5348) );
  AND2X1 U6584 ( .A(\RF[14][49] ), .B(n10729), .Y(n1268) );
  INVX1 U6585 ( .A(n1268), .Y(n5349) );
  AND2X1 U6586 ( .A(\RF[15][50] ), .B(n10731), .Y(n1203) );
  INVX1 U6587 ( .A(n1203), .Y(n5350) );
  AND2X1 U6588 ( .A(\RF[16][45] ), .B(n10733), .Y(n1133) );
  INVX1 U6589 ( .A(n1133), .Y(n5351) );
  AND2X1 U6590 ( .A(\RF[16][32] ), .B(n10733), .Y(n1120) );
  INVX1 U6591 ( .A(n1120), .Y(n5352) );
  AND2X1 U6592 ( .A(\RF[16][13] ), .B(n10734), .Y(n1101) );
  INVX1 U6593 ( .A(n1101), .Y(n5353) );
  AND2X1 U6594 ( .A(\RF[16][1] ), .B(n10733), .Y(n1089) );
  INVX1 U6595 ( .A(n1089), .Y(n5354) );
  AND2X1 U6596 ( .A(\RF[16][0] ), .B(n10733), .Y(n1088) );
  INVX1 U6597 ( .A(n1088), .Y(n5355) );
  AND2X1 U6598 ( .A(\RF[17][37] ), .B(n10735), .Y(n1060) );
  INVX1 U6599 ( .A(n1060), .Y(n5356) );
  AND2X1 U6600 ( .A(\RF[17][26] ), .B(n10736), .Y(n1049) );
  INVX1 U6601 ( .A(n1049), .Y(n5357) );
  AND2X1 U6602 ( .A(\RF[17][14] ), .B(n10735), .Y(n1037) );
  INVX1 U6603 ( .A(n1037), .Y(n5358) );
  AND2X1 U6604 ( .A(\RF[17][2] ), .B(n10736), .Y(n1025) );
  INVX1 U6605 ( .A(n1025), .Y(n5359) );
  AND2X1 U6606 ( .A(\RF[18][39] ), .B(n10737), .Y(n997) );
  INVX1 U6607 ( .A(n997), .Y(n5360) );
  AND2X1 U6608 ( .A(\RF[18][27] ), .B(n10738), .Y(n985) );
  INVX1 U6609 ( .A(n985), .Y(n5361) );
  AND2X1 U6610 ( .A(\RF[18][15] ), .B(n10737), .Y(n973) );
  INVX1 U6611 ( .A(n973), .Y(n5362) );
  AND2X1 U6612 ( .A(\RF[18][3] ), .B(n10738), .Y(n961) );
  INVX1 U6613 ( .A(n961), .Y(n5363) );
  AND2X1 U6614 ( .A(\RF[19][40] ), .B(n10739), .Y(n933) );
  INVX1 U6615 ( .A(n933), .Y(n5364) );
  AND2X1 U6616 ( .A(\RF[19][28] ), .B(n10740), .Y(n921) );
  INVX1 U6617 ( .A(n921), .Y(n5365) );
  AND2X1 U6618 ( .A(\RF[19][16] ), .B(n10739), .Y(n909) );
  INVX1 U6619 ( .A(n909), .Y(n5366) );
  AND2X1 U6620 ( .A(\RF[19][4] ), .B(n10740), .Y(n897) );
  INVX1 U6621 ( .A(n897), .Y(n5367) );
  AND2X1 U6622 ( .A(\RF[20][41] ), .B(n10741), .Y(n869) );
  INVX1 U6623 ( .A(n869), .Y(n5368) );
  AND2X1 U6624 ( .A(\RF[20][29] ), .B(n10742), .Y(n857) );
  INVX1 U6625 ( .A(n857), .Y(n5369) );
  AND2X1 U6626 ( .A(\RF[20][17] ), .B(n10741), .Y(n845) );
  INVX1 U6627 ( .A(n845), .Y(n5370) );
  AND2X1 U6628 ( .A(\RF[20][5] ), .B(n10742), .Y(n833) );
  INVX1 U6629 ( .A(n833), .Y(n5371) );
  AND2X1 U6630 ( .A(\RF[21][38] ), .B(n10744), .Y(n801) );
  INVX1 U6631 ( .A(n801), .Y(n5372) );
  AND2X1 U6632 ( .A(\RF[21][30] ), .B(n10743), .Y(n793) );
  INVX1 U6633 ( .A(n793), .Y(n5373) );
  AND2X1 U6634 ( .A(\RF[21][18] ), .B(n10743), .Y(n781) );
  INVX1 U6635 ( .A(n781), .Y(n5374) );
  AND2X1 U6636 ( .A(\RF[21][6] ), .B(n10744), .Y(n769) );
  INVX1 U6637 ( .A(n769), .Y(n5375) );
  AND2X1 U6638 ( .A(\RF[22][43] ), .B(n10745), .Y(n741) );
  INVX1 U6639 ( .A(n741), .Y(n5376) );
  AND2X1 U6640 ( .A(\RF[22][31] ), .B(n10746), .Y(n729) );
  INVX1 U6641 ( .A(n729), .Y(n5377) );
  AND2X1 U6642 ( .A(\RF[22][19] ), .B(n10745), .Y(n717) );
  INVX1 U6643 ( .A(n717), .Y(n5378) );
  AND2X1 U6644 ( .A(\RF[22][7] ), .B(n10746), .Y(n705) );
  INVX1 U6645 ( .A(n705), .Y(n5379) );
  AND2X1 U6646 ( .A(\RF[23][47] ), .B(n10747), .Y(n679) );
  INVX1 U6647 ( .A(n679), .Y(n5380) );
  AND2X1 U6648 ( .A(\RF[23][25] ), .B(n10747), .Y(n657) );
  INVX1 U6649 ( .A(n657), .Y(n5381) );
  AND2X1 U6650 ( .A(\RF[23][20] ), .B(n10748), .Y(n652) );
  INVX1 U6651 ( .A(n652), .Y(n5382) );
  AND2X1 U6652 ( .A(\RF[23][8] ), .B(n10748), .Y(n640) );
  INVX1 U6653 ( .A(n640), .Y(n5383) );
  AND2X1 U6654 ( .A(\RF[24][45] ), .B(n10749), .Y(n610) );
  INVX1 U6655 ( .A(n610), .Y(n5384) );
  AND2X1 U6656 ( .A(\RF[24][32] ), .B(n10749), .Y(n597) );
  INVX1 U6657 ( .A(n597), .Y(n5385) );
  AND2X1 U6658 ( .A(\RF[24][13] ), .B(n10750), .Y(n578) );
  INVX1 U6659 ( .A(n578), .Y(n5386) );
  AND2X1 U6660 ( .A(\RF[24][1] ), .B(n10749), .Y(n566) );
  INVX1 U6661 ( .A(n566), .Y(n5387) );
  AND2X1 U6662 ( .A(\RF[24][0] ), .B(n10749), .Y(n565) );
  INVX1 U6663 ( .A(n565), .Y(n5388) );
  AND2X1 U6664 ( .A(\RF[25][37] ), .B(n10751), .Y(n536) );
  INVX1 U6665 ( .A(n536), .Y(n5389) );
  AND2X1 U6666 ( .A(\RF[25][26] ), .B(n10752), .Y(n525) );
  INVX1 U6667 ( .A(n525), .Y(n5390) );
  AND2X1 U6668 ( .A(\RF[25][14] ), .B(n10751), .Y(n513) );
  INVX1 U6669 ( .A(n513), .Y(n5391) );
  AND2X1 U6670 ( .A(\RF[25][2] ), .B(n10752), .Y(n501) );
  INVX1 U6671 ( .A(n501), .Y(n5392) );
  AND2X1 U6672 ( .A(\RF[26][39] ), .B(n10753), .Y(n472) );
  INVX1 U6673 ( .A(n472), .Y(n5393) );
  AND2X1 U6674 ( .A(\RF[26][27] ), .B(n10754), .Y(n460) );
  INVX1 U6675 ( .A(n460), .Y(n5394) );
  AND2X1 U6676 ( .A(\RF[26][15] ), .B(n10753), .Y(n448) );
  INVX1 U6677 ( .A(n448), .Y(n5395) );
  AND2X1 U6678 ( .A(\RF[26][3] ), .B(n10754), .Y(n436) );
  INVX1 U6679 ( .A(n436), .Y(n5396) );
  AND2X1 U6680 ( .A(\RF[27][40] ), .B(n10755), .Y(n407) );
  INVX1 U6681 ( .A(n407), .Y(n5397) );
  AND2X1 U6682 ( .A(\RF[27][28] ), .B(n10756), .Y(n395) );
  INVX1 U6683 ( .A(n395), .Y(n5398) );
  AND2X1 U6684 ( .A(\RF[27][16] ), .B(n10755), .Y(n383) );
  INVX1 U6685 ( .A(n383), .Y(n5399) );
  AND2X1 U6686 ( .A(\RF[27][4] ), .B(n10756), .Y(n371) );
  INVX1 U6687 ( .A(n371), .Y(n5400) );
  AND2X1 U6688 ( .A(\RF[28][41] ), .B(n10757), .Y(n342) );
  INVX1 U6689 ( .A(n342), .Y(n5401) );
  AND2X1 U6690 ( .A(\RF[28][29] ), .B(n10758), .Y(n330) );
  INVX1 U6691 ( .A(n330), .Y(n5402) );
  AND2X1 U6692 ( .A(\RF[28][17] ), .B(n10757), .Y(n318) );
  INVX1 U6693 ( .A(n318), .Y(n5403) );
  AND2X1 U6694 ( .A(\RF[28][5] ), .B(n10758), .Y(n306) );
  INVX1 U6695 ( .A(n306), .Y(n5404) );
  AND2X1 U6696 ( .A(\RF[29][38] ), .B(n10760), .Y(n273) );
  INVX1 U6697 ( .A(n273), .Y(n5405) );
  AND2X1 U6698 ( .A(\RF[29][30] ), .B(n10759), .Y(n265) );
  INVX1 U6699 ( .A(n265), .Y(n5406) );
  AND2X1 U6700 ( .A(\RF[29][18] ), .B(n10759), .Y(n253) );
  INVX1 U6701 ( .A(n253), .Y(n5407) );
  AND2X1 U6702 ( .A(\RF[29][6] ), .B(n10760), .Y(n241) );
  INVX1 U6703 ( .A(n241), .Y(n5408) );
  AND2X1 U6704 ( .A(\RF[30][43] ), .B(n10761), .Y(n212) );
  INVX1 U6705 ( .A(n212), .Y(n5409) );
  AND2X1 U6706 ( .A(\RF[30][31] ), .B(n10762), .Y(n200) );
  INVX1 U6707 ( .A(n200), .Y(n5410) );
  AND2X1 U6708 ( .A(\RF[30][19] ), .B(n10761), .Y(n188) );
  INVX1 U6709 ( .A(n188), .Y(n5411) );
  AND2X1 U6710 ( .A(\RF[30][7] ), .B(n10762), .Y(n176) );
  INVX1 U6711 ( .A(n176), .Y(n5412) );
  AND2X1 U6712 ( .A(\RF[31][47] ), .B(n10763), .Y(n133) );
  INVX1 U6713 ( .A(n133), .Y(n5413) );
  AND2X1 U6714 ( .A(\RF[31][25] ), .B(n10763), .Y(n89) );
  INVX1 U6715 ( .A(n89), .Y(n5414) );
  AND2X1 U6716 ( .A(\RF[31][20] ), .B(n10764), .Y(n79) );
  INVX1 U6717 ( .A(n79), .Y(n5415) );
  AND2X1 U6718 ( .A(\RF[31][8] ), .B(n10764), .Y(n55) );
  INVX1 U6719 ( .A(n55), .Y(n5416) );
  BUFX2 U6720 ( .A(n564), .Y(n5417) );
  AND2X1 U6721 ( .A(\RF[0][58] ), .B(n10702), .Y(n2188) );
  INVX1 U6722 ( .A(n2188), .Y(n5418) );
  AND2X1 U6723 ( .A(\RF[0][48] ), .B(n10702), .Y(n2178) );
  INVX1 U6724 ( .A(n2178), .Y(n5419) );
  AND2X1 U6725 ( .A(\RF[1][57] ), .B(n10704), .Y(n2122) );
  INVX1 U6726 ( .A(n2122), .Y(n5420) );
  AND2X1 U6727 ( .A(\RF[1][46] ), .B(n10704), .Y(n2111) );
  INVX1 U6728 ( .A(n2111), .Y(n5421) );
  AND2X1 U6729 ( .A(\RF[1][24] ), .B(n10703), .Y(n2089) );
  INVX1 U6730 ( .A(n2089), .Y(n5422) );
  AND2X1 U6731 ( .A(\RF[2][50] ), .B(n10706), .Y(n2050) );
  INVX1 U6732 ( .A(n2050), .Y(n5423) );
  AND2X1 U6733 ( .A(\RF[3][61] ), .B(n10708), .Y(n1996) );
  INVX1 U6734 ( .A(n1996), .Y(n5424) );
  AND2X1 U6735 ( .A(\RF[3][53] ), .B(n10708), .Y(n1988) );
  INVX1 U6736 ( .A(n1988), .Y(n5425) );
  AND2X1 U6737 ( .A(\RF[3][49] ), .B(n10708), .Y(n1984) );
  INVX1 U6738 ( .A(n1984), .Y(n5426) );
  AND2X1 U6739 ( .A(\RF[4][37] ), .B(n10710), .Y(n1907) );
  INVX1 U6740 ( .A(n1907), .Y(n5427) );
  AND2X1 U6741 ( .A(\RF[4][26] ), .B(n10710), .Y(n1896) );
  INVX1 U6742 ( .A(n1896), .Y(n5428) );
  AND2X1 U6743 ( .A(\RF[4][14] ), .B(n10710), .Y(n1884) );
  INVX1 U6744 ( .A(n1884), .Y(n5429) );
  AND2X1 U6745 ( .A(\RF[4][2] ), .B(n10710), .Y(n1872) );
  INVX1 U6746 ( .A(n1872), .Y(n5430) );
  AND2X1 U6747 ( .A(\RF[5][45] ), .B(n10712), .Y(n1850) );
  INVX1 U6748 ( .A(n1850), .Y(n5431) );
  AND2X1 U6749 ( .A(\RF[5][32] ), .B(n10712), .Y(n1837) );
  INVX1 U6750 ( .A(n1837), .Y(n5432) );
  AND2X1 U6751 ( .A(\RF[5][13] ), .B(n10712), .Y(n1818) );
  INVX1 U6752 ( .A(n1818), .Y(n5433) );
  AND2X1 U6753 ( .A(\RF[5][1] ), .B(n10712), .Y(n1806) );
  INVX1 U6754 ( .A(n1806), .Y(n5434) );
  AND2X1 U6755 ( .A(\RF[5][0] ), .B(n10711), .Y(n1805) );
  INVX1 U6756 ( .A(n1805), .Y(n5435) );
  AND2X1 U6757 ( .A(\RF[6][40] ), .B(n10714), .Y(n1780) );
  INVX1 U6758 ( .A(n1780), .Y(n5436) );
  AND2X1 U6759 ( .A(\RF[6][28] ), .B(n10714), .Y(n1768) );
  INVX1 U6760 ( .A(n1768), .Y(n5437) );
  AND2X1 U6761 ( .A(\RF[6][16] ), .B(n10714), .Y(n1756) );
  INVX1 U6762 ( .A(n1756), .Y(n5438) );
  AND2X1 U6763 ( .A(\RF[6][4] ), .B(n10714), .Y(n1744) );
  INVX1 U6764 ( .A(n1744), .Y(n5439) );
  AND2X1 U6765 ( .A(\RF[7][39] ), .B(n10716), .Y(n1713) );
  INVX1 U6766 ( .A(n1713), .Y(n5440) );
  AND2X1 U6767 ( .A(\RF[7][27] ), .B(n10716), .Y(n1701) );
  INVX1 U6768 ( .A(n1701), .Y(n5441) );
  AND2X1 U6769 ( .A(\RF[7][15] ), .B(n10716), .Y(n1689) );
  INVX1 U6770 ( .A(n1689), .Y(n5442) );
  AND2X1 U6771 ( .A(\RF[7][3] ), .B(n10716), .Y(n1677) );
  INVX1 U6772 ( .A(n1677), .Y(n5443) );
  AND2X1 U6773 ( .A(\RF[8][38] ), .B(n10718), .Y(n1647) );
  INVX1 U6774 ( .A(n1647), .Y(n5444) );
  AND2X1 U6775 ( .A(\RF[8][30] ), .B(n10718), .Y(n1639) );
  INVX1 U6776 ( .A(n1639), .Y(n5445) );
  AND2X1 U6777 ( .A(\RF[8][18] ), .B(n10718), .Y(n1627) );
  INVX1 U6778 ( .A(n1627), .Y(n5446) );
  AND2X1 U6779 ( .A(\RF[8][6] ), .B(n10718), .Y(n1615) );
  INVX1 U6780 ( .A(n1615), .Y(n5447) );
  AND2X1 U6781 ( .A(\RF[9][41] ), .B(n10720), .Y(n1585) );
  INVX1 U6782 ( .A(n1585), .Y(n5448) );
  AND2X1 U6783 ( .A(\RF[9][29] ), .B(n10720), .Y(n1573) );
  INVX1 U6784 ( .A(n1573), .Y(n5449) );
  AND2X1 U6785 ( .A(\RF[9][17] ), .B(n10720), .Y(n1561) );
  INVX1 U6786 ( .A(n1561), .Y(n5450) );
  AND2X1 U6787 ( .A(\RF[9][5] ), .B(n10720), .Y(n1549) );
  INVX1 U6788 ( .A(n1549), .Y(n5451) );
  AND2X1 U6789 ( .A(\RF[10][47] ), .B(n10722), .Y(n1526) );
  INVX1 U6790 ( .A(n1526), .Y(n5452) );
  AND2X1 U6791 ( .A(\RF[10][25] ), .B(n10722), .Y(n1504) );
  INVX1 U6792 ( .A(n1504), .Y(n5453) );
  AND2X1 U6793 ( .A(\RF[10][20] ), .B(n10722), .Y(n1499) );
  INVX1 U6794 ( .A(n1499), .Y(n5454) );
  AND2X1 U6795 ( .A(\RF[10][8] ), .B(n10722), .Y(n1487) );
  INVX1 U6796 ( .A(n1487), .Y(n5455) );
  AND2X1 U6797 ( .A(\RF[11][43] ), .B(n10724), .Y(n1457) );
  INVX1 U6798 ( .A(n1457), .Y(n5456) );
  AND2X1 U6799 ( .A(\RF[11][31] ), .B(n10724), .Y(n1445) );
  INVX1 U6800 ( .A(n1445), .Y(n5457) );
  AND2X1 U6801 ( .A(\RF[11][19] ), .B(n10724), .Y(n1433) );
  INVX1 U6802 ( .A(n1433), .Y(n5458) );
  AND2X1 U6803 ( .A(\RF[11][7] ), .B(n10724), .Y(n1421) );
  INVX1 U6804 ( .A(n1421), .Y(n5459) );
  AND2X1 U6805 ( .A(\RF[12][58] ), .B(n10726), .Y(n1407) );
  INVX1 U6806 ( .A(n1407), .Y(n5460) );
  AND2X1 U6807 ( .A(\RF[12][48] ), .B(n10726), .Y(n1397) );
  INVX1 U6808 ( .A(n1397), .Y(n5461) );
  AND2X1 U6809 ( .A(\RF[13][57] ), .B(n10728), .Y(n1341) );
  INVX1 U6810 ( .A(n1341), .Y(n5462) );
  AND2X1 U6811 ( .A(\RF[13][46] ), .B(n10728), .Y(n1330) );
  INVX1 U6812 ( .A(n1330), .Y(n5463) );
  AND2X1 U6813 ( .A(\RF[13][24] ), .B(n10727), .Y(n1308) );
  INVX1 U6814 ( .A(n1308), .Y(n5464) );
  AND2X1 U6815 ( .A(\RF[14][50] ), .B(n10730), .Y(n1269) );
  INVX1 U6816 ( .A(n1269), .Y(n5465) );
  AND2X1 U6817 ( .A(\RF[15][61] ), .B(n10732), .Y(n1214) );
  INVX1 U6818 ( .A(n1214), .Y(n5466) );
  AND2X1 U6819 ( .A(\RF[15][53] ), .B(n10732), .Y(n1206) );
  INVX1 U6820 ( .A(n1206), .Y(n5467) );
  AND2X1 U6821 ( .A(\RF[15][49] ), .B(n10732), .Y(n1202) );
  INVX1 U6822 ( .A(n1202), .Y(n5468) );
  AND2X1 U6823 ( .A(\RF[16][37] ), .B(n10734), .Y(n1125) );
  INVX1 U6824 ( .A(n1125), .Y(n5469) );
  AND2X1 U6825 ( .A(\RF[16][26] ), .B(n10734), .Y(n1114) );
  INVX1 U6826 ( .A(n1114), .Y(n5470) );
  AND2X1 U6827 ( .A(\RF[16][14] ), .B(n10734), .Y(n1102) );
  INVX1 U6828 ( .A(n1102), .Y(n5471) );
  AND2X1 U6829 ( .A(\RF[16][2] ), .B(n10734), .Y(n1090) );
  INVX1 U6830 ( .A(n1090), .Y(n5472) );
  AND2X1 U6831 ( .A(\RF[17][45] ), .B(n10736), .Y(n1068) );
  INVX1 U6832 ( .A(n1068), .Y(n5473) );
  AND2X1 U6833 ( .A(\RF[17][32] ), .B(n10736), .Y(n1055) );
  INVX1 U6834 ( .A(n1055), .Y(n5474) );
  AND2X1 U6835 ( .A(\RF[17][13] ), .B(n10736), .Y(n1036) );
  INVX1 U6836 ( .A(n1036), .Y(n5475) );
  AND2X1 U6837 ( .A(\RF[17][1] ), .B(n10736), .Y(n1024) );
  INVX1 U6838 ( .A(n1024), .Y(n5476) );
  AND2X1 U6839 ( .A(\RF[17][0] ), .B(n10735), .Y(n1023) );
  INVX1 U6840 ( .A(n1023), .Y(n5477) );
  AND2X1 U6841 ( .A(\RF[18][40] ), .B(n10738), .Y(n998) );
  INVX1 U6842 ( .A(n998), .Y(n5478) );
  AND2X1 U6843 ( .A(\RF[18][28] ), .B(n10738), .Y(n986) );
  INVX1 U6844 ( .A(n986), .Y(n5479) );
  AND2X1 U6845 ( .A(\RF[18][16] ), .B(n10738), .Y(n974) );
  INVX1 U6846 ( .A(n974), .Y(n5480) );
  AND2X1 U6847 ( .A(\RF[18][4] ), .B(n10738), .Y(n962) );
  INVX1 U6848 ( .A(n962), .Y(n5481) );
  AND2X1 U6849 ( .A(\RF[19][39] ), .B(n10740), .Y(n932) );
  INVX1 U6850 ( .A(n932), .Y(n5482) );
  AND2X1 U6851 ( .A(\RF[19][27] ), .B(n10740), .Y(n920) );
  INVX1 U6852 ( .A(n920), .Y(n5483) );
  AND2X1 U6853 ( .A(\RF[19][15] ), .B(n10740), .Y(n908) );
  INVX1 U6854 ( .A(n908), .Y(n5484) );
  AND2X1 U6855 ( .A(\RF[19][3] ), .B(n10740), .Y(n896) );
  INVX1 U6856 ( .A(n896), .Y(n5485) );
  AND2X1 U6857 ( .A(\RF[20][38] ), .B(n10742), .Y(n866) );
  INVX1 U6858 ( .A(n866), .Y(n5486) );
  AND2X1 U6859 ( .A(\RF[20][30] ), .B(n10742), .Y(n858) );
  INVX1 U6860 ( .A(n858), .Y(n5487) );
  AND2X1 U6861 ( .A(\RF[20][18] ), .B(n10742), .Y(n846) );
  INVX1 U6862 ( .A(n846), .Y(n5488) );
  AND2X1 U6863 ( .A(\RF[20][6] ), .B(n10742), .Y(n834) );
  INVX1 U6864 ( .A(n834), .Y(n5489) );
  AND2X1 U6865 ( .A(\RF[21][41] ), .B(n10744), .Y(n804) );
  INVX1 U6866 ( .A(n804), .Y(n5490) );
  AND2X1 U6867 ( .A(\RF[21][29] ), .B(n10744), .Y(n792) );
  INVX1 U6868 ( .A(n792), .Y(n5491) );
  AND2X1 U6869 ( .A(\RF[21][17] ), .B(n10744), .Y(n780) );
  INVX1 U6870 ( .A(n780), .Y(n5492) );
  AND2X1 U6871 ( .A(\RF[21][5] ), .B(n10744), .Y(n768) );
  INVX1 U6872 ( .A(n768), .Y(n5493) );
  AND2X1 U6873 ( .A(\RF[22][47] ), .B(n10746), .Y(n745) );
  INVX1 U6874 ( .A(n745), .Y(n5494) );
  AND2X1 U6875 ( .A(\RF[22][25] ), .B(n10746), .Y(n723) );
  INVX1 U6876 ( .A(n723), .Y(n5495) );
  AND2X1 U6877 ( .A(\RF[22][20] ), .B(n10746), .Y(n718) );
  INVX1 U6878 ( .A(n718), .Y(n5496) );
  AND2X1 U6879 ( .A(\RF[22][8] ), .B(n10746), .Y(n706) );
  INVX1 U6880 ( .A(n706), .Y(n5497) );
  AND2X1 U6881 ( .A(\RF[23][43] ), .B(n10748), .Y(n675) );
  INVX1 U6882 ( .A(n675), .Y(n5498) );
  AND2X1 U6883 ( .A(\RF[23][31] ), .B(n10748), .Y(n663) );
  INVX1 U6884 ( .A(n663), .Y(n5499) );
  AND2X1 U6885 ( .A(\RF[23][19] ), .B(n10748), .Y(n651) );
  INVX1 U6886 ( .A(n651), .Y(n5500) );
  AND2X1 U6887 ( .A(\RF[23][7] ), .B(n10748), .Y(n639) );
  INVX1 U6888 ( .A(n639), .Y(n5501) );
  AND2X1 U6889 ( .A(\RF[24][37] ), .B(n10750), .Y(n602) );
  INVX1 U6890 ( .A(n602), .Y(n5502) );
  AND2X1 U6891 ( .A(\RF[24][26] ), .B(n10750), .Y(n591) );
  INVX1 U6892 ( .A(n591), .Y(n5503) );
  AND2X1 U6893 ( .A(\RF[24][14] ), .B(n10750), .Y(n579) );
  INVX1 U6894 ( .A(n579), .Y(n5504) );
  AND2X1 U6895 ( .A(\RF[24][2] ), .B(n10750), .Y(n567) );
  INVX1 U6896 ( .A(n567), .Y(n5505) );
  AND2X1 U6897 ( .A(\RF[25][45] ), .B(n10752), .Y(n544) );
  INVX1 U6898 ( .A(n544), .Y(n5506) );
  AND2X1 U6899 ( .A(\RF[25][32] ), .B(n10752), .Y(n531) );
  INVX1 U6900 ( .A(n531), .Y(n5507) );
  AND2X1 U6901 ( .A(\RF[25][13] ), .B(n10752), .Y(n512) );
  INVX1 U6902 ( .A(n512), .Y(n5508) );
  AND2X1 U6903 ( .A(\RF[25][1] ), .B(n10752), .Y(n500) );
  INVX1 U6904 ( .A(n500), .Y(n5509) );
  AND2X1 U6905 ( .A(\RF[25][0] ), .B(n10751), .Y(n499) );
  INVX1 U6906 ( .A(n499), .Y(n5510) );
  AND2X1 U6907 ( .A(\RF[26][40] ), .B(n10754), .Y(n473) );
  INVX1 U6908 ( .A(n473), .Y(n5511) );
  AND2X1 U6909 ( .A(\RF[26][28] ), .B(n10754), .Y(n461) );
  INVX1 U6910 ( .A(n461), .Y(n5512) );
  AND2X1 U6911 ( .A(\RF[26][16] ), .B(n10754), .Y(n449) );
  INVX1 U6912 ( .A(n449), .Y(n5513) );
  AND2X1 U6913 ( .A(\RF[26][4] ), .B(n10754), .Y(n437) );
  INVX1 U6914 ( .A(n437), .Y(n5514) );
  AND2X1 U6915 ( .A(\RF[27][39] ), .B(n10756), .Y(n406) );
  INVX1 U6916 ( .A(n406), .Y(n5515) );
  AND2X1 U6917 ( .A(\RF[27][27] ), .B(n10756), .Y(n394) );
  INVX1 U6918 ( .A(n394), .Y(n5516) );
  AND2X1 U6919 ( .A(\RF[27][15] ), .B(n10756), .Y(n382) );
  INVX1 U6920 ( .A(n382), .Y(n5517) );
  AND2X1 U6921 ( .A(\RF[27][3] ), .B(n10756), .Y(n370) );
  INVX1 U6922 ( .A(n370), .Y(n5518) );
  AND2X1 U6923 ( .A(\RF[28][38] ), .B(n10758), .Y(n339) );
  INVX1 U6924 ( .A(n339), .Y(n5519) );
  AND2X1 U6925 ( .A(\RF[28][30] ), .B(n10758), .Y(n331) );
  INVX1 U6926 ( .A(n331), .Y(n5520) );
  AND2X1 U6927 ( .A(\RF[28][18] ), .B(n10758), .Y(n319) );
  INVX1 U6928 ( .A(n319), .Y(n5521) );
  AND2X1 U6929 ( .A(\RF[28][6] ), .B(n10758), .Y(n307) );
  INVX1 U6930 ( .A(n307), .Y(n5522) );
  AND2X1 U6931 ( .A(\RF[29][41] ), .B(n10760), .Y(n276) );
  INVX1 U6932 ( .A(n276), .Y(n5523) );
  AND2X1 U6933 ( .A(\RF[29][29] ), .B(n10760), .Y(n264) );
  INVX1 U6934 ( .A(n264), .Y(n5524) );
  AND2X1 U6935 ( .A(\RF[29][17] ), .B(n10760), .Y(n252) );
  INVX1 U6936 ( .A(n252), .Y(n5525) );
  AND2X1 U6937 ( .A(\RF[29][5] ), .B(n10760), .Y(n240) );
  INVX1 U6938 ( .A(n240), .Y(n5526) );
  AND2X1 U6939 ( .A(\RF[30][47] ), .B(n10762), .Y(n216) );
  INVX1 U6940 ( .A(n216), .Y(n5527) );
  AND2X1 U6941 ( .A(\RF[30][25] ), .B(n10762), .Y(n194) );
  INVX1 U6942 ( .A(n194), .Y(n5528) );
  AND2X1 U6943 ( .A(\RF[30][20] ), .B(n10762), .Y(n189) );
  INVX1 U6944 ( .A(n189), .Y(n5529) );
  AND2X1 U6945 ( .A(\RF[30][8] ), .B(n10762), .Y(n177) );
  INVX1 U6946 ( .A(n177), .Y(n5530) );
  AND2X1 U6947 ( .A(\RF[31][43] ), .B(n10764), .Y(n125) );
  INVX1 U6948 ( .A(n125), .Y(n5531) );
  AND2X1 U6949 ( .A(\RF[31][31] ), .B(n10764), .Y(n101) );
  INVX1 U6950 ( .A(n101), .Y(n5532) );
  AND2X1 U6951 ( .A(\RF[31][19] ), .B(n10764), .Y(n77) );
  INVX1 U6952 ( .A(n77), .Y(n5533) );
  AND2X1 U6953 ( .A(\RF[31][7] ), .B(n10764), .Y(n53) );
  INVX1 U6954 ( .A(n53), .Y(n5534) );
  BUFX2 U6955 ( .A(n498), .Y(n5535) );
  AND2X1 U6956 ( .A(\RF[0][61] ), .B(n10702), .Y(n2191) );
  INVX1 U6957 ( .A(n2191), .Y(n5536) );
  AND2X1 U6958 ( .A(\RF[0][53] ), .B(n10701), .Y(n2183) );
  INVX1 U6959 ( .A(n2183), .Y(n5537) );
  AND2X1 U6960 ( .A(\RF[0][49] ), .B(n10701), .Y(n2179) );
  INVX1 U6961 ( .A(n2179), .Y(n5538) );
  AND2X1 U6962 ( .A(\RF[1][50] ), .B(n10703), .Y(n2115) );
  INVX1 U6963 ( .A(n2115), .Y(n5539) );
  AND2X1 U6964 ( .A(\RF[2][57] ), .B(n10705), .Y(n2057) );
  INVX1 U6965 ( .A(n2057), .Y(n5540) );
  AND2X1 U6966 ( .A(\RF[2][46] ), .B(n10706), .Y(n2046) );
  INVX1 U6967 ( .A(n2046), .Y(n5541) );
  AND2X1 U6968 ( .A(\RF[2][24] ), .B(n10705), .Y(n2024) );
  INVX1 U6969 ( .A(n2024), .Y(n5542) );
  AND2X1 U6970 ( .A(\RF[3][58] ), .B(n10707), .Y(n1993) );
  INVX1 U6971 ( .A(n1993), .Y(n5543) );
  AND2X1 U6972 ( .A(\RF[3][48] ), .B(n10707), .Y(n1983) );
  INVX1 U6973 ( .A(n1983), .Y(n5544) );
  AND2X1 U6974 ( .A(\RF[4][39] ), .B(n10709), .Y(n1909) );
  INVX1 U6975 ( .A(n1909), .Y(n5545) );
  AND2X1 U6976 ( .A(\RF[4][27] ), .B(n10709), .Y(n1897) );
  INVX1 U6977 ( .A(n1897), .Y(n5546) );
  AND2X1 U6978 ( .A(\RF[4][15] ), .B(n10710), .Y(n1885) );
  INVX1 U6979 ( .A(n1885), .Y(n5547) );
  AND2X1 U6980 ( .A(\RF[4][3] ), .B(n10709), .Y(n1873) );
  INVX1 U6981 ( .A(n1873), .Y(n5548) );
  AND2X1 U6982 ( .A(\RF[5][40] ), .B(n10711), .Y(n1845) );
  INVX1 U6983 ( .A(n1845), .Y(n5549) );
  AND2X1 U6984 ( .A(\RF[5][28] ), .B(n10712), .Y(n1833) );
  INVX1 U6985 ( .A(n1833), .Y(n5550) );
  AND2X1 U6986 ( .A(\RF[5][16] ), .B(n10711), .Y(n1821) );
  INVX1 U6987 ( .A(n1821), .Y(n5551) );
  AND2X1 U6988 ( .A(\RF[5][4] ), .B(n10711), .Y(n1809) );
  INVX1 U6989 ( .A(n1809), .Y(n5552) );
  AND2X1 U6990 ( .A(\RF[6][45] ), .B(n10714), .Y(n1785) );
  INVX1 U6991 ( .A(n1785), .Y(n5553) );
  AND2X1 U6992 ( .A(\RF[6][32] ), .B(n10713), .Y(n1772) );
  INVX1 U6993 ( .A(n1772), .Y(n5554) );
  AND2X1 U6994 ( .A(\RF[6][13] ), .B(n10713), .Y(n1753) );
  INVX1 U6995 ( .A(n1753), .Y(n5555) );
  AND2X1 U6996 ( .A(\RF[6][1] ), .B(n10713), .Y(n1741) );
  INVX1 U6997 ( .A(n1741), .Y(n5556) );
  AND2X1 U6998 ( .A(\RF[6][0] ), .B(n10713), .Y(n1740) );
  INVX1 U6999 ( .A(n1740), .Y(n5557) );
  AND2X1 U7000 ( .A(\RF[7][37] ), .B(n10715), .Y(n1711) );
  INVX1 U7001 ( .A(n1711), .Y(n5558) );
  AND2X1 U7002 ( .A(\RF[7][26] ), .B(n10716), .Y(n1700) );
  INVX1 U7003 ( .A(n1700), .Y(n5559) );
  AND2X1 U7004 ( .A(\RF[7][14] ), .B(n10715), .Y(n1688) );
  INVX1 U7005 ( .A(n1688), .Y(n5560) );
  AND2X1 U7006 ( .A(\RF[7][2] ), .B(n10715), .Y(n1676) );
  INVX1 U7007 ( .A(n1676), .Y(n5561) );
  AND2X1 U7008 ( .A(\RF[8][43] ), .B(n10717), .Y(n1652) );
  INVX1 U7009 ( .A(n1652), .Y(n5562) );
  AND2X1 U7010 ( .A(\RF[8][31] ), .B(n10718), .Y(n1640) );
  INVX1 U7011 ( .A(n1640), .Y(n5563) );
  AND2X1 U7012 ( .A(\RF[8][19] ), .B(n10717), .Y(n1628) );
  INVX1 U7013 ( .A(n1628), .Y(n5564) );
  AND2X1 U7014 ( .A(\RF[8][7] ), .B(n10717), .Y(n1616) );
  INVX1 U7015 ( .A(n1616), .Y(n5565) );
  AND2X1 U7016 ( .A(\RF[9][47] ), .B(n10719), .Y(n1591) );
  INVX1 U7017 ( .A(n1591), .Y(n5566) );
  AND2X1 U7018 ( .A(\RF[9][25] ), .B(n10719), .Y(n1569) );
  INVX1 U7019 ( .A(n1569), .Y(n5567) );
  AND2X1 U7020 ( .A(\RF[9][20] ), .B(n10720), .Y(n1564) );
  INVX1 U7021 ( .A(n1564), .Y(n5568) );
  AND2X1 U7022 ( .A(\RF[9][8] ), .B(n10719), .Y(n1552) );
  INVX1 U7023 ( .A(n1552), .Y(n5569) );
  AND2X1 U7024 ( .A(\RF[10][41] ), .B(n10721), .Y(n1520) );
  INVX1 U7025 ( .A(n1520), .Y(n5570) );
  AND2X1 U7026 ( .A(\RF[10][29] ), .B(n10722), .Y(n1508) );
  INVX1 U7027 ( .A(n1508), .Y(n5571) );
  AND2X1 U7028 ( .A(\RF[10][17] ), .B(n10721), .Y(n1496) );
  INVX1 U7029 ( .A(n1496), .Y(n5572) );
  AND2X1 U7030 ( .A(\RF[10][5] ), .B(n10721), .Y(n1484) );
  INVX1 U7031 ( .A(n1484), .Y(n5573) );
  AND2X1 U7032 ( .A(\RF[11][38] ), .B(n10724), .Y(n1452) );
  INVX1 U7033 ( .A(n1452), .Y(n5574) );
  AND2X1 U7034 ( .A(\RF[11][30] ), .B(n10723), .Y(n1444) );
  INVX1 U7035 ( .A(n1444), .Y(n5575) );
  AND2X1 U7036 ( .A(\RF[11][18] ), .B(n10723), .Y(n1432) );
  INVX1 U7037 ( .A(n1432), .Y(n5576) );
  AND2X1 U7038 ( .A(\RF[11][6] ), .B(n10723), .Y(n1420) );
  INVX1 U7039 ( .A(n1420), .Y(n5577) );
  AND2X1 U7040 ( .A(\RF[12][61] ), .B(n10726), .Y(n1410) );
  INVX1 U7041 ( .A(n1410), .Y(n5578) );
  AND2X1 U7042 ( .A(\RF[12][53] ), .B(n10725), .Y(n1402) );
  INVX1 U7043 ( .A(n1402), .Y(n5579) );
  AND2X1 U7044 ( .A(\RF[12][49] ), .B(n10725), .Y(n1398) );
  INVX1 U7045 ( .A(n1398), .Y(n5580) );
  AND2X1 U7046 ( .A(\RF[13][50] ), .B(n10727), .Y(n1334) );
  INVX1 U7047 ( .A(n1334), .Y(n5581) );
  AND2X1 U7048 ( .A(\RF[14][57] ), .B(n10729), .Y(n1276) );
  INVX1 U7049 ( .A(n1276), .Y(n5582) );
  AND2X1 U7050 ( .A(\RF[14][46] ), .B(n10730), .Y(n1265) );
  INVX1 U7051 ( .A(n1265), .Y(n5583) );
  AND2X1 U7052 ( .A(\RF[14][24] ), .B(n10729), .Y(n1243) );
  INVX1 U7053 ( .A(n1243), .Y(n5584) );
  AND2X1 U7054 ( .A(\RF[15][58] ), .B(n10731), .Y(n1211) );
  INVX1 U7055 ( .A(n1211), .Y(n5585) );
  AND2X1 U7056 ( .A(\RF[15][48] ), .B(n10731), .Y(n1201) );
  INVX1 U7057 ( .A(n1201), .Y(n5586) );
  AND2X1 U7058 ( .A(\RF[16][39] ), .B(n10733), .Y(n1127) );
  INVX1 U7059 ( .A(n1127), .Y(n5587) );
  AND2X1 U7060 ( .A(\RF[16][27] ), .B(n10733), .Y(n1115) );
  INVX1 U7061 ( .A(n1115), .Y(n5588) );
  AND2X1 U7062 ( .A(\RF[16][15] ), .B(n10734), .Y(n1103) );
  INVX1 U7063 ( .A(n1103), .Y(n5589) );
  AND2X1 U7064 ( .A(\RF[16][3] ), .B(n10733), .Y(n1091) );
  INVX1 U7065 ( .A(n1091), .Y(n5590) );
  AND2X1 U7066 ( .A(\RF[17][40] ), .B(n10735), .Y(n1063) );
  INVX1 U7067 ( .A(n1063), .Y(n5591) );
  AND2X1 U7068 ( .A(\RF[17][28] ), .B(n10736), .Y(n1051) );
  INVX1 U7069 ( .A(n1051), .Y(n5592) );
  AND2X1 U7070 ( .A(\RF[17][16] ), .B(n10735), .Y(n1039) );
  INVX1 U7071 ( .A(n1039), .Y(n5593) );
  AND2X1 U7072 ( .A(\RF[17][4] ), .B(n10735), .Y(n1027) );
  INVX1 U7073 ( .A(n1027), .Y(n5594) );
  AND2X1 U7074 ( .A(\RF[18][45] ), .B(n10738), .Y(n1003) );
  INVX1 U7075 ( .A(n1003), .Y(n5595) );
  AND2X1 U7076 ( .A(\RF[18][32] ), .B(n10737), .Y(n990) );
  INVX1 U7077 ( .A(n990), .Y(n5596) );
  AND2X1 U7078 ( .A(\RF[18][13] ), .B(n10737), .Y(n971) );
  INVX1 U7079 ( .A(n971), .Y(n5597) );
  AND2X1 U7080 ( .A(\RF[18][1] ), .B(n10737), .Y(n959) );
  INVX1 U7081 ( .A(n959), .Y(n5598) );
  AND2X1 U7082 ( .A(\RF[18][0] ), .B(n10737), .Y(n958) );
  INVX1 U7083 ( .A(n958), .Y(n5599) );
  AND2X1 U7084 ( .A(\RF[19][37] ), .B(n10739), .Y(n930) );
  INVX1 U7085 ( .A(n930), .Y(n5600) );
  AND2X1 U7086 ( .A(\RF[19][26] ), .B(n10740), .Y(n919) );
  INVX1 U7087 ( .A(n919), .Y(n5601) );
  AND2X1 U7088 ( .A(\RF[19][14] ), .B(n10739), .Y(n907) );
  INVX1 U7089 ( .A(n907), .Y(n5602) );
  AND2X1 U7090 ( .A(\RF[19][2] ), .B(n10739), .Y(n895) );
  INVX1 U7091 ( .A(n895), .Y(n5603) );
  AND2X1 U7092 ( .A(\RF[20][43] ), .B(n10741), .Y(n871) );
  INVX1 U7093 ( .A(n871), .Y(n5604) );
  AND2X1 U7094 ( .A(\RF[20][31] ), .B(n10742), .Y(n859) );
  INVX1 U7095 ( .A(n859), .Y(n5605) );
  AND2X1 U7096 ( .A(\RF[20][19] ), .B(n10741), .Y(n847) );
  INVX1 U7097 ( .A(n847), .Y(n5606) );
  AND2X1 U7098 ( .A(\RF[20][7] ), .B(n10741), .Y(n835) );
  INVX1 U7099 ( .A(n835), .Y(n5607) );
  AND2X1 U7100 ( .A(\RF[21][47] ), .B(n10743), .Y(n810) );
  INVX1 U7101 ( .A(n810), .Y(n5608) );
  AND2X1 U7102 ( .A(\RF[21][25] ), .B(n10743), .Y(n788) );
  INVX1 U7103 ( .A(n788), .Y(n5609) );
  AND2X1 U7104 ( .A(\RF[21][20] ), .B(n10744), .Y(n783) );
  INVX1 U7105 ( .A(n783), .Y(n5610) );
  AND2X1 U7106 ( .A(\RF[21][8] ), .B(n10743), .Y(n771) );
  INVX1 U7107 ( .A(n771), .Y(n5611) );
  AND2X1 U7108 ( .A(\RF[22][41] ), .B(n10745), .Y(n739) );
  INVX1 U7109 ( .A(n739), .Y(n5612) );
  AND2X1 U7110 ( .A(\RF[22][29] ), .B(n10746), .Y(n727) );
  INVX1 U7111 ( .A(n727), .Y(n5613) );
  AND2X1 U7112 ( .A(\RF[22][17] ), .B(n10745), .Y(n715) );
  INVX1 U7113 ( .A(n715), .Y(n5614) );
  AND2X1 U7114 ( .A(\RF[22][5] ), .B(n10745), .Y(n703) );
  INVX1 U7115 ( .A(n703), .Y(n5615) );
  AND2X1 U7116 ( .A(\RF[23][38] ), .B(n10748), .Y(n670) );
  INVX1 U7117 ( .A(n670), .Y(n5616) );
  AND2X1 U7118 ( .A(\RF[23][30] ), .B(n10747), .Y(n662) );
  INVX1 U7119 ( .A(n662), .Y(n5617) );
  AND2X1 U7120 ( .A(\RF[23][18] ), .B(n10747), .Y(n650) );
  INVX1 U7121 ( .A(n650), .Y(n5618) );
  AND2X1 U7122 ( .A(\RF[23][6] ), .B(n10747), .Y(n638) );
  INVX1 U7123 ( .A(n638), .Y(n5619) );
  AND2X1 U7124 ( .A(\RF[24][39] ), .B(n10749), .Y(n604) );
  INVX1 U7125 ( .A(n604), .Y(n5620) );
  AND2X1 U7126 ( .A(\RF[24][27] ), .B(n10749), .Y(n592) );
  INVX1 U7127 ( .A(n592), .Y(n5621) );
  AND2X1 U7128 ( .A(\RF[24][15] ), .B(n10750), .Y(n580) );
  INVX1 U7129 ( .A(n580), .Y(n5622) );
  AND2X1 U7130 ( .A(\RF[24][3] ), .B(n10749), .Y(n568) );
  INVX1 U7131 ( .A(n568), .Y(n5623) );
  AND2X1 U7132 ( .A(\RF[25][40] ), .B(n10751), .Y(n539) );
  INVX1 U7133 ( .A(n539), .Y(n5624) );
  AND2X1 U7134 ( .A(\RF[25][28] ), .B(n10752), .Y(n527) );
  INVX1 U7135 ( .A(n527), .Y(n5625) );
  AND2X1 U7136 ( .A(\RF[25][16] ), .B(n10751), .Y(n515) );
  INVX1 U7137 ( .A(n515), .Y(n5626) );
  AND2X1 U7138 ( .A(\RF[25][4] ), .B(n10751), .Y(n503) );
  INVX1 U7139 ( .A(n503), .Y(n5627) );
  AND2X1 U7140 ( .A(\RF[26][45] ), .B(n10754), .Y(n478) );
  INVX1 U7141 ( .A(n478), .Y(n5628) );
  AND2X1 U7142 ( .A(\RF[26][32] ), .B(n10753), .Y(n465) );
  INVX1 U7143 ( .A(n465), .Y(n5629) );
  AND2X1 U7144 ( .A(\RF[26][13] ), .B(n10753), .Y(n446) );
  INVX1 U7145 ( .A(n446), .Y(n5630) );
  AND2X1 U7146 ( .A(\RF[26][1] ), .B(n10753), .Y(n434) );
  INVX1 U7147 ( .A(n434), .Y(n5631) );
  AND2X1 U7148 ( .A(\RF[26][0] ), .B(n10753), .Y(n433) );
  INVX1 U7149 ( .A(n433), .Y(n5632) );
  AND2X1 U7150 ( .A(\RF[27][37] ), .B(n10755), .Y(n404) );
  INVX1 U7151 ( .A(n404), .Y(n5633) );
  AND2X1 U7152 ( .A(\RF[27][26] ), .B(n10756), .Y(n393) );
  INVX1 U7153 ( .A(n393), .Y(n5634) );
  AND2X1 U7154 ( .A(\RF[27][14] ), .B(n10755), .Y(n381) );
  INVX1 U7155 ( .A(n381), .Y(n5635) );
  AND2X1 U7156 ( .A(\RF[27][2] ), .B(n10755), .Y(n369) );
  INVX1 U7157 ( .A(n369), .Y(n5636) );
  AND2X1 U7158 ( .A(\RF[28][43] ), .B(n10757), .Y(n344) );
  INVX1 U7159 ( .A(n344), .Y(n5637) );
  AND2X1 U7160 ( .A(\RF[28][31] ), .B(n10758), .Y(n332) );
  INVX1 U7161 ( .A(n332), .Y(n5638) );
  AND2X1 U7162 ( .A(\RF[28][19] ), .B(n10757), .Y(n320) );
  INVX1 U7163 ( .A(n320), .Y(n5639) );
  AND2X1 U7164 ( .A(\RF[28][7] ), .B(n10757), .Y(n308) );
  INVX1 U7165 ( .A(n308), .Y(n5640) );
  AND2X1 U7166 ( .A(\RF[29][47] ), .B(n10759), .Y(n282) );
  INVX1 U7167 ( .A(n282), .Y(n5641) );
  AND2X1 U7168 ( .A(\RF[29][25] ), .B(n10759), .Y(n260) );
  INVX1 U7169 ( .A(n260), .Y(n5642) );
  AND2X1 U7170 ( .A(\RF[29][20] ), .B(n10760), .Y(n255) );
  INVX1 U7171 ( .A(n255), .Y(n5643) );
  AND2X1 U7172 ( .A(\RF[29][8] ), .B(n10759), .Y(n243) );
  INVX1 U7173 ( .A(n243), .Y(n5644) );
  AND2X1 U7174 ( .A(\RF[30][41] ), .B(n10761), .Y(n210) );
  INVX1 U7175 ( .A(n210), .Y(n5645) );
  AND2X1 U7176 ( .A(\RF[30][29] ), .B(n10762), .Y(n198) );
  INVX1 U7177 ( .A(n198), .Y(n5646) );
  AND2X1 U7178 ( .A(\RF[30][17] ), .B(n10761), .Y(n186) );
  INVX1 U7179 ( .A(n186), .Y(n5647) );
  AND2X1 U7180 ( .A(\RF[30][5] ), .B(n10761), .Y(n174) );
  INVX1 U7181 ( .A(n174), .Y(n5648) );
  AND2X1 U7182 ( .A(\RF[31][38] ), .B(n10764), .Y(n115) );
  INVX1 U7183 ( .A(n115), .Y(n5649) );
  AND2X1 U7184 ( .A(\RF[31][30] ), .B(n10763), .Y(n99) );
  INVX1 U7185 ( .A(n99), .Y(n5650) );
  AND2X1 U7186 ( .A(\RF[31][18] ), .B(n10763), .Y(n75) );
  INVX1 U7187 ( .A(n75), .Y(n5651) );
  AND2X1 U7188 ( .A(\RF[31][6] ), .B(n10763), .Y(n51) );
  INVX1 U7189 ( .A(n51), .Y(n5652) );
  BUFX2 U7190 ( .A(n366), .Y(n5653) );
  AND2X1 U7191 ( .A(\RF[0][50] ), .B(n10701), .Y(n2180) );
  INVX1 U7192 ( .A(n2180), .Y(n5654) );
  AND2X1 U7193 ( .A(\RF[1][61] ), .B(n10704), .Y(n2126) );
  INVX1 U7194 ( .A(n2126), .Y(n5655) );
  AND2X1 U7195 ( .A(\RF[1][53] ), .B(n10703), .Y(n2118) );
  INVX1 U7196 ( .A(n2118), .Y(n5656) );
  AND2X1 U7197 ( .A(\RF[1][49] ), .B(n10703), .Y(n2114) );
  INVX1 U7198 ( .A(n2114), .Y(n5657) );
  AND2X1 U7199 ( .A(\RF[2][58] ), .B(n10705), .Y(n2058) );
  INVX1 U7200 ( .A(n2058), .Y(n5658) );
  AND2X1 U7201 ( .A(\RF[2][48] ), .B(n10706), .Y(n2048) );
  INVX1 U7202 ( .A(n2048), .Y(n5659) );
  AND2X1 U7203 ( .A(\RF[3][57] ), .B(n10707), .Y(n1992) );
  INVX1 U7204 ( .A(n1992), .Y(n5660) );
  AND2X1 U7205 ( .A(\RF[3][46] ), .B(n10707), .Y(n1981) );
  INVX1 U7206 ( .A(n1981), .Y(n5661) );
  AND2X1 U7207 ( .A(\RF[3][24] ), .B(n10708), .Y(n1959) );
  INVX1 U7208 ( .A(n1959), .Y(n5662) );
  AND2X1 U7209 ( .A(\RF[4][40] ), .B(n10710), .Y(n1910) );
  INVX1 U7210 ( .A(n1910), .Y(n5663) );
  AND2X1 U7211 ( .A(\RF[4][28] ), .B(n10709), .Y(n1898) );
  INVX1 U7212 ( .A(n1898), .Y(n5664) );
  AND2X1 U7213 ( .A(\RF[4][16] ), .B(n10710), .Y(n1886) );
  INVX1 U7214 ( .A(n1886), .Y(n5665) );
  AND2X1 U7215 ( .A(\RF[4][4] ), .B(n10709), .Y(n1874) );
  INVX1 U7216 ( .A(n1874), .Y(n5666) );
  AND2X1 U7217 ( .A(\RF[5][39] ), .B(n10712), .Y(n1844) );
  INVX1 U7218 ( .A(n1844), .Y(n5667) );
  AND2X1 U7219 ( .A(\RF[5][27] ), .B(n10712), .Y(n1832) );
  INVX1 U7220 ( .A(n1832), .Y(n5668) );
  AND2X1 U7221 ( .A(\RF[5][15] ), .B(n10711), .Y(n1820) );
  INVX1 U7222 ( .A(n1820), .Y(n5669) );
  AND2X1 U7223 ( .A(\RF[5][3] ), .B(n10711), .Y(n1808) );
  INVX1 U7224 ( .A(n1808), .Y(n5670) );
  AND2X1 U7225 ( .A(\RF[6][37] ), .B(n10714), .Y(n1777) );
  INVX1 U7226 ( .A(n1777), .Y(n5671) );
  AND2X1 U7227 ( .A(\RF[6][26] ), .B(n10714), .Y(n1766) );
  INVX1 U7228 ( .A(n1766), .Y(n5672) );
  AND2X1 U7229 ( .A(\RF[6][14] ), .B(n10713), .Y(n1754) );
  INVX1 U7230 ( .A(n1754), .Y(n5673) );
  AND2X1 U7231 ( .A(\RF[6][2] ), .B(n10713), .Y(n1742) );
  INVX1 U7232 ( .A(n1742), .Y(n5674) );
  AND2X1 U7233 ( .A(\RF[7][45] ), .B(n10716), .Y(n1719) );
  INVX1 U7234 ( .A(n1719), .Y(n5675) );
  AND2X1 U7235 ( .A(\RF[7][32] ), .B(n10716), .Y(n1706) );
  INVX1 U7236 ( .A(n1706), .Y(n5676) );
  AND2X1 U7237 ( .A(\RF[7][13] ), .B(n10715), .Y(n1687) );
  INVX1 U7238 ( .A(n1687), .Y(n5677) );
  AND2X1 U7239 ( .A(\RF[7][1] ), .B(n10715), .Y(n1675) );
  INVX1 U7240 ( .A(n1675), .Y(n5678) );
  AND2X1 U7241 ( .A(\RF[7][0] ), .B(n10715), .Y(n1674) );
  INVX1 U7242 ( .A(n1674), .Y(n5679) );
  AND2X1 U7243 ( .A(\RF[8][47] ), .B(n10718), .Y(n1656) );
  INVX1 U7244 ( .A(n1656), .Y(n5680) );
  AND2X1 U7245 ( .A(\RF[8][25] ), .B(n10717), .Y(n1634) );
  INVX1 U7246 ( .A(n1634), .Y(n5681) );
  AND2X1 U7247 ( .A(\RF[8][20] ), .B(n10718), .Y(n1629) );
  INVX1 U7248 ( .A(n1629), .Y(n5682) );
  AND2X1 U7249 ( .A(\RF[8][8] ), .B(n10717), .Y(n1617) );
  INVX1 U7250 ( .A(n1617), .Y(n5683) );
  AND2X1 U7251 ( .A(\RF[9][43] ), .B(n10720), .Y(n1587) );
  INVX1 U7252 ( .A(n1587), .Y(n5684) );
  AND2X1 U7253 ( .A(\RF[9][31] ), .B(n10720), .Y(n1575) );
  INVX1 U7254 ( .A(n1575), .Y(n5685) );
  AND2X1 U7255 ( .A(\RF[9][19] ), .B(n10719), .Y(n1563) );
  INVX1 U7256 ( .A(n1563), .Y(n5686) );
  AND2X1 U7257 ( .A(\RF[9][7] ), .B(n10719), .Y(n1551) );
  INVX1 U7258 ( .A(n1551), .Y(n5687) );
  AND2X1 U7259 ( .A(\RF[10][38] ), .B(n10722), .Y(n1517) );
  INVX1 U7260 ( .A(n1517), .Y(n5688) );
  AND2X1 U7261 ( .A(\RF[10][30] ), .B(n10722), .Y(n1509) );
  INVX1 U7262 ( .A(n1509), .Y(n5689) );
  AND2X1 U7263 ( .A(\RF[10][18] ), .B(n10721), .Y(n1497) );
  INVX1 U7264 ( .A(n1497), .Y(n5690) );
  AND2X1 U7265 ( .A(\RF[10][6] ), .B(n10721), .Y(n1485) );
  INVX1 U7266 ( .A(n1485), .Y(n5691) );
  AND2X1 U7267 ( .A(\RF[11][41] ), .B(n10724), .Y(n1455) );
  INVX1 U7268 ( .A(n1455), .Y(n5692) );
  AND2X1 U7269 ( .A(\RF[11][29] ), .B(n10724), .Y(n1443) );
  INVX1 U7270 ( .A(n1443), .Y(n5693) );
  AND2X1 U7271 ( .A(\RF[11][17] ), .B(n10723), .Y(n1431) );
  INVX1 U7272 ( .A(n1431), .Y(n5694) );
  AND2X1 U7273 ( .A(\RF[11][5] ), .B(n10723), .Y(n1419) );
  INVX1 U7274 ( .A(n1419), .Y(n5695) );
  AND2X1 U7275 ( .A(\RF[12][50] ), .B(n10725), .Y(n1399) );
  INVX1 U7276 ( .A(n1399), .Y(n5696) );
  AND2X1 U7277 ( .A(\RF[13][61] ), .B(n10728), .Y(n1345) );
  INVX1 U7278 ( .A(n1345), .Y(n5697) );
  AND2X1 U7279 ( .A(\RF[13][53] ), .B(n10727), .Y(n1337) );
  INVX1 U7280 ( .A(n1337), .Y(n5698) );
  AND2X1 U7281 ( .A(\RF[13][49] ), .B(n10727), .Y(n1333) );
  INVX1 U7282 ( .A(n1333), .Y(n5699) );
  AND2X1 U7283 ( .A(\RF[14][58] ), .B(n10729), .Y(n1277) );
  INVX1 U7284 ( .A(n1277), .Y(n5700) );
  AND2X1 U7285 ( .A(\RF[14][48] ), .B(n10730), .Y(n1267) );
  INVX1 U7286 ( .A(n1267), .Y(n5701) );
  AND2X1 U7287 ( .A(\RF[15][57] ), .B(n10731), .Y(n1210) );
  INVX1 U7288 ( .A(n1210), .Y(n5702) );
  AND2X1 U7289 ( .A(\RF[15][46] ), .B(n10731), .Y(n1199) );
  INVX1 U7290 ( .A(n1199), .Y(n5703) );
  AND2X1 U7291 ( .A(\RF[15][24] ), .B(n10732), .Y(n1177) );
  INVX1 U7292 ( .A(n1177), .Y(n5704) );
  AND2X1 U7293 ( .A(\RF[16][40] ), .B(n10734), .Y(n1128) );
  INVX1 U7294 ( .A(n1128), .Y(n5705) );
  AND2X1 U7295 ( .A(\RF[16][28] ), .B(n10733), .Y(n1116) );
  INVX1 U7296 ( .A(n1116), .Y(n5706) );
  AND2X1 U7297 ( .A(\RF[16][16] ), .B(n10734), .Y(n1104) );
  INVX1 U7298 ( .A(n1104), .Y(n5707) );
  AND2X1 U7299 ( .A(\RF[16][4] ), .B(n10733), .Y(n1092) );
  INVX1 U7300 ( .A(n1092), .Y(n5708) );
  AND2X1 U7301 ( .A(\RF[17][39] ), .B(n10736), .Y(n1062) );
  INVX1 U7302 ( .A(n1062), .Y(n5709) );
  AND2X1 U7303 ( .A(\RF[17][27] ), .B(n10736), .Y(n1050) );
  INVX1 U7304 ( .A(n1050), .Y(n5710) );
  AND2X1 U7305 ( .A(\RF[17][15] ), .B(n10735), .Y(n1038) );
  INVX1 U7306 ( .A(n1038), .Y(n5711) );
  AND2X1 U7307 ( .A(\RF[17][3] ), .B(n10735), .Y(n1026) );
  INVX1 U7308 ( .A(n1026), .Y(n5712) );
  AND2X1 U7309 ( .A(\RF[18][37] ), .B(n10738), .Y(n995) );
  INVX1 U7310 ( .A(n995), .Y(n5713) );
  AND2X1 U7311 ( .A(\RF[18][26] ), .B(n10738), .Y(n984) );
  INVX1 U7312 ( .A(n984), .Y(n5714) );
  AND2X1 U7313 ( .A(\RF[18][14] ), .B(n10737), .Y(n972) );
  INVX1 U7314 ( .A(n972), .Y(n5715) );
  AND2X1 U7315 ( .A(\RF[18][2] ), .B(n10737), .Y(n960) );
  INVX1 U7316 ( .A(n960), .Y(n5716) );
  AND2X1 U7317 ( .A(\RF[19][45] ), .B(n10740), .Y(n938) );
  INVX1 U7318 ( .A(n938), .Y(n5717) );
  AND2X1 U7319 ( .A(\RF[19][32] ), .B(n10740), .Y(n925) );
  INVX1 U7320 ( .A(n925), .Y(n5718) );
  AND2X1 U7321 ( .A(\RF[19][13] ), .B(n10739), .Y(n906) );
  INVX1 U7322 ( .A(n906), .Y(n5719) );
  AND2X1 U7323 ( .A(\RF[19][1] ), .B(n10739), .Y(n894) );
  INVX1 U7324 ( .A(n894), .Y(n5720) );
  AND2X1 U7325 ( .A(\RF[19][0] ), .B(n10739), .Y(n893) );
  INVX1 U7326 ( .A(n893), .Y(n5721) );
  AND2X1 U7327 ( .A(\RF[20][47] ), .B(n10742), .Y(n875) );
  INVX1 U7328 ( .A(n875), .Y(n5722) );
  AND2X1 U7329 ( .A(\RF[20][25] ), .B(n10741), .Y(n853) );
  INVX1 U7330 ( .A(n853), .Y(n5723) );
  AND2X1 U7331 ( .A(\RF[20][20] ), .B(n10742), .Y(n848) );
  INVX1 U7332 ( .A(n848), .Y(n5724) );
  AND2X1 U7333 ( .A(\RF[20][8] ), .B(n10741), .Y(n836) );
  INVX1 U7334 ( .A(n836), .Y(n5725) );
  AND2X1 U7335 ( .A(\RF[21][43] ), .B(n10744), .Y(n806) );
  INVX1 U7336 ( .A(n806), .Y(n5726) );
  AND2X1 U7337 ( .A(\RF[21][31] ), .B(n10744), .Y(n794) );
  INVX1 U7338 ( .A(n794), .Y(n5727) );
  AND2X1 U7339 ( .A(\RF[21][19] ), .B(n10743), .Y(n782) );
  INVX1 U7340 ( .A(n782), .Y(n5728) );
  AND2X1 U7341 ( .A(\RF[21][7] ), .B(n10743), .Y(n770) );
  INVX1 U7342 ( .A(n770), .Y(n5729) );
  AND2X1 U7343 ( .A(\RF[22][38] ), .B(n10746), .Y(n736) );
  INVX1 U7344 ( .A(n736), .Y(n5730) );
  AND2X1 U7345 ( .A(\RF[22][30] ), .B(n10746), .Y(n728) );
  INVX1 U7346 ( .A(n728), .Y(n5731) );
  AND2X1 U7347 ( .A(\RF[22][18] ), .B(n10745), .Y(n716) );
  INVX1 U7348 ( .A(n716), .Y(n5732) );
  AND2X1 U7349 ( .A(\RF[22][6] ), .B(n10745), .Y(n704) );
  INVX1 U7350 ( .A(n704), .Y(n5733) );
  AND2X1 U7351 ( .A(\RF[23][41] ), .B(n10748), .Y(n673) );
  INVX1 U7352 ( .A(n673), .Y(n5734) );
  AND2X1 U7353 ( .A(\RF[23][29] ), .B(n10748), .Y(n661) );
  INVX1 U7354 ( .A(n661), .Y(n5735) );
  AND2X1 U7355 ( .A(\RF[23][17] ), .B(n10747), .Y(n649) );
  INVX1 U7356 ( .A(n649), .Y(n5736) );
  AND2X1 U7357 ( .A(\RF[23][5] ), .B(n10747), .Y(n637) );
  INVX1 U7358 ( .A(n637), .Y(n5737) );
  AND2X1 U7359 ( .A(\RF[24][40] ), .B(n10750), .Y(n605) );
  INVX1 U7360 ( .A(n605), .Y(n5738) );
  AND2X1 U7361 ( .A(\RF[24][28] ), .B(n10749), .Y(n593) );
  INVX1 U7362 ( .A(n593), .Y(n5739) );
  AND2X1 U7363 ( .A(\RF[24][16] ), .B(n10750), .Y(n581) );
  INVX1 U7364 ( .A(n581), .Y(n5740) );
  AND2X1 U7365 ( .A(\RF[24][4] ), .B(n10749), .Y(n569) );
  INVX1 U7366 ( .A(n569), .Y(n5741) );
  AND2X1 U7367 ( .A(\RF[25][39] ), .B(n10752), .Y(n538) );
  INVX1 U7368 ( .A(n538), .Y(n5742) );
  AND2X1 U7369 ( .A(\RF[25][27] ), .B(n10752), .Y(n526) );
  INVX1 U7370 ( .A(n526), .Y(n5743) );
  AND2X1 U7371 ( .A(\RF[25][15] ), .B(n10751), .Y(n514) );
  INVX1 U7372 ( .A(n514), .Y(n5744) );
  AND2X1 U7373 ( .A(\RF[25][3] ), .B(n10751), .Y(n502) );
  INVX1 U7374 ( .A(n502), .Y(n5745) );
  AND2X1 U7375 ( .A(\RF[26][37] ), .B(n10754), .Y(n470) );
  INVX1 U7376 ( .A(n470), .Y(n5746) );
  AND2X1 U7377 ( .A(\RF[26][26] ), .B(n10754), .Y(n459) );
  INVX1 U7378 ( .A(n459), .Y(n5747) );
  AND2X1 U7379 ( .A(\RF[26][14] ), .B(n10753), .Y(n447) );
  INVX1 U7380 ( .A(n447), .Y(n5748) );
  AND2X1 U7381 ( .A(\RF[26][2] ), .B(n10753), .Y(n435) );
  INVX1 U7382 ( .A(n435), .Y(n5749) );
  AND2X1 U7383 ( .A(\RF[27][45] ), .B(n10756), .Y(n412) );
  INVX1 U7384 ( .A(n412), .Y(n5750) );
  AND2X1 U7385 ( .A(\RF[27][32] ), .B(n10756), .Y(n399) );
  INVX1 U7386 ( .A(n399), .Y(n5751) );
  AND2X1 U7387 ( .A(\RF[27][13] ), .B(n10755), .Y(n380) );
  INVX1 U7388 ( .A(n380), .Y(n5752) );
  AND2X1 U7389 ( .A(\RF[27][1] ), .B(n10755), .Y(n368) );
  INVX1 U7390 ( .A(n368), .Y(n5753) );
  AND2X1 U7391 ( .A(\RF[27][0] ), .B(n10755), .Y(n367) );
  INVX1 U7392 ( .A(n367), .Y(n5754) );
  AND2X1 U7393 ( .A(\RF[28][47] ), .B(n10758), .Y(n348) );
  INVX1 U7394 ( .A(n348), .Y(n5755) );
  AND2X1 U7395 ( .A(\RF[28][25] ), .B(n10757), .Y(n326) );
  INVX1 U7396 ( .A(n326), .Y(n5756) );
  AND2X1 U7397 ( .A(\RF[28][20] ), .B(n10758), .Y(n321) );
  INVX1 U7398 ( .A(n321), .Y(n5757) );
  AND2X1 U7399 ( .A(\RF[28][8] ), .B(n10757), .Y(n309) );
  INVX1 U7400 ( .A(n309), .Y(n5758) );
  AND2X1 U7401 ( .A(\RF[29][43] ), .B(n10760), .Y(n278) );
  INVX1 U7402 ( .A(n278), .Y(n5759) );
  AND2X1 U7403 ( .A(\RF[29][31] ), .B(n10760), .Y(n266) );
  INVX1 U7404 ( .A(n266), .Y(n5760) );
  AND2X1 U7405 ( .A(\RF[29][19] ), .B(n10759), .Y(n254) );
  INVX1 U7406 ( .A(n254), .Y(n5761) );
  AND2X1 U7407 ( .A(\RF[29][7] ), .B(n10759), .Y(n242) );
  INVX1 U7408 ( .A(n242), .Y(n5762) );
  AND2X1 U7409 ( .A(\RF[30][38] ), .B(n10762), .Y(n207) );
  INVX1 U7410 ( .A(n207), .Y(n5763) );
  AND2X1 U7411 ( .A(\RF[30][30] ), .B(n10762), .Y(n199) );
  INVX1 U7412 ( .A(n199), .Y(n5764) );
  AND2X1 U7413 ( .A(\RF[30][18] ), .B(n10761), .Y(n187) );
  INVX1 U7414 ( .A(n187), .Y(n5765) );
  AND2X1 U7415 ( .A(\RF[30][6] ), .B(n10761), .Y(n175) );
  INVX1 U7416 ( .A(n175), .Y(n5766) );
  AND2X1 U7417 ( .A(\RF[31][41] ), .B(n10764), .Y(n121) );
  INVX1 U7418 ( .A(n121), .Y(n5767) );
  AND2X1 U7419 ( .A(\RF[31][29] ), .B(n10764), .Y(n97) );
  INVX1 U7420 ( .A(n97), .Y(n5768) );
  AND2X1 U7421 ( .A(\RF[31][17] ), .B(n10763), .Y(n73) );
  INVX1 U7422 ( .A(n73), .Y(n5769) );
  AND2X1 U7423 ( .A(\RF[31][5] ), .B(n10763), .Y(n49) );
  INVX1 U7424 ( .A(n49), .Y(n5770) );
  BUFX2 U7425 ( .A(n432), .Y(n5771) );
  BUFX2 U7426 ( .A(n300), .Y(n5772) );
  BUFX2 U7427 ( .A(n234), .Y(n5773) );
  BUFX2 U7428 ( .A(n168), .Y(n5774) );
  AND2X1 U7429 ( .A(\RF[0][44] ), .B(n10701), .Y(n2174) );
  INVX1 U7430 ( .A(n2174), .Y(n5775) );
  AND2X1 U7431 ( .A(\RF[0][33] ), .B(n10702), .Y(n2163) );
  INVX1 U7432 ( .A(n2163), .Y(n5776) );
  AND2X1 U7433 ( .A(\RF[0][21] ), .B(n10702), .Y(n2151) );
  INVX1 U7434 ( .A(n2151), .Y(n5777) );
  AND2X1 U7435 ( .A(\RF[0][9] ), .B(n10702), .Y(n2139) );
  INVX1 U7436 ( .A(n2139), .Y(n5778) );
  AND2X1 U7437 ( .A(\RF[1][63] ), .B(n10703), .Y(n2128) );
  INVX1 U7438 ( .A(n2128), .Y(n5779) );
  AND2X1 U7439 ( .A(\RF[1][34] ), .B(n10704), .Y(n2099) );
  INVX1 U7440 ( .A(n2099), .Y(n5780) );
  AND2X1 U7441 ( .A(\RF[1][22] ), .B(n10703), .Y(n2087) );
  INVX1 U7442 ( .A(n2087), .Y(n5781) );
  AND2X1 U7443 ( .A(\RF[1][10] ), .B(n10704), .Y(n2075) );
  INVX1 U7444 ( .A(n2075), .Y(n5782) );
  AND2X1 U7445 ( .A(\RF[2][56] ), .B(n10706), .Y(n2056) );
  INVX1 U7446 ( .A(n2056), .Y(n5783) );
  AND2X1 U7447 ( .A(\RF[2][35] ), .B(n10706), .Y(n2035) );
  INVX1 U7448 ( .A(n2035), .Y(n5784) );
  AND2X1 U7449 ( .A(\RF[2][23] ), .B(n10706), .Y(n2023) );
  INVX1 U7450 ( .A(n2023), .Y(n5785) );
  AND2X1 U7451 ( .A(\RF[2][11] ), .B(n10706), .Y(n2011) );
  INVX1 U7452 ( .A(n2011), .Y(n5786) );
  AND2X1 U7453 ( .A(\RF[3][59] ), .B(n10707), .Y(n1994) );
  INVX1 U7454 ( .A(n1994), .Y(n5787) );
  AND2X1 U7455 ( .A(\RF[3][42] ), .B(n10708), .Y(n1977) );
  INVX1 U7456 ( .A(n1977), .Y(n5788) );
  AND2X1 U7457 ( .A(\RF[3][36] ), .B(n10708), .Y(n1971) );
  INVX1 U7458 ( .A(n1971), .Y(n5789) );
  AND2X1 U7459 ( .A(\RF[3][12] ), .B(n10708), .Y(n1947) );
  INVX1 U7460 ( .A(n1947), .Y(n5790) );
  AND2X1 U7461 ( .A(\RF[4][41] ), .B(n10709), .Y(n1911) );
  INVX1 U7462 ( .A(n1911), .Y(n5791) );
  AND2X1 U7463 ( .A(\RF[4][29] ), .B(n10710), .Y(n1899) );
  INVX1 U7464 ( .A(n1899), .Y(n5792) );
  AND2X1 U7465 ( .A(\RF[4][17] ), .B(n10710), .Y(n1887) );
  INVX1 U7466 ( .A(n1887), .Y(n5793) );
  AND2X1 U7467 ( .A(\RF[4][5] ), .B(n10709), .Y(n1875) );
  INVX1 U7468 ( .A(n1875), .Y(n5794) );
  AND2X1 U7469 ( .A(\RF[5][38] ), .B(n10712), .Y(n1843) );
  INVX1 U7470 ( .A(n1843), .Y(n5795) );
  AND2X1 U7471 ( .A(\RF[5][30] ), .B(n10711), .Y(n1835) );
  INVX1 U7472 ( .A(n1835), .Y(n5796) );
  AND2X1 U7473 ( .A(\RF[5][18] ), .B(n10712), .Y(n1823) );
  INVX1 U7474 ( .A(n1823), .Y(n5797) );
  AND2X1 U7475 ( .A(\RF[5][6] ), .B(n10712), .Y(n1811) );
  INVX1 U7476 ( .A(n1811), .Y(n5798) );
  AND2X1 U7477 ( .A(\RF[6][43] ), .B(n10713), .Y(n1783) );
  INVX1 U7478 ( .A(n1783), .Y(n5799) );
  AND2X1 U7479 ( .A(\RF[6][31] ), .B(n10714), .Y(n1771) );
  INVX1 U7480 ( .A(n1771), .Y(n5800) );
  AND2X1 U7481 ( .A(\RF[6][19] ), .B(n10714), .Y(n1759) );
  INVX1 U7482 ( .A(n1759), .Y(n5801) );
  AND2X1 U7483 ( .A(\RF[6][7] ), .B(n10714), .Y(n1747) );
  INVX1 U7484 ( .A(n1747), .Y(n5802) );
  AND2X1 U7485 ( .A(\RF[7][47] ), .B(n10715), .Y(n1721) );
  INVX1 U7486 ( .A(n1721), .Y(n5803) );
  AND2X1 U7487 ( .A(\RF[7][25] ), .B(n10716), .Y(n1699) );
  INVX1 U7488 ( .A(n1699), .Y(n5804) );
  AND2X1 U7489 ( .A(\RF[7][20] ), .B(n10716), .Y(n1694) );
  INVX1 U7490 ( .A(n1694), .Y(n5805) );
  AND2X1 U7491 ( .A(\RF[7][8] ), .B(n10716), .Y(n1682) );
  INVX1 U7492 ( .A(n1682), .Y(n5806) );
  AND2X1 U7493 ( .A(\RF[8][45] ), .B(n10718), .Y(n1654) );
  INVX1 U7494 ( .A(n1654), .Y(n5807) );
  AND2X1 U7495 ( .A(\RF[8][32] ), .B(n10717), .Y(n1641) );
  INVX1 U7496 ( .A(n1641), .Y(n5808) );
  AND2X1 U7497 ( .A(\RF[8][13] ), .B(n10718), .Y(n1622) );
  INVX1 U7498 ( .A(n1622), .Y(n5809) );
  AND2X1 U7499 ( .A(\RF[8][1] ), .B(n10718), .Y(n1610) );
  INVX1 U7500 ( .A(n1610), .Y(n5810) );
  AND2X1 U7501 ( .A(\RF[8][0] ), .B(n10717), .Y(n1609) );
  INVX1 U7502 ( .A(n1609), .Y(n5811) );
  AND2X1 U7503 ( .A(\RF[9][37] ), .B(n10719), .Y(n1581) );
  INVX1 U7504 ( .A(n1581), .Y(n5812) );
  AND2X1 U7505 ( .A(\RF[9][26] ), .B(n10720), .Y(n1570) );
  INVX1 U7506 ( .A(n1570), .Y(n5813) );
  AND2X1 U7507 ( .A(\RF[9][14] ), .B(n10720), .Y(n1558) );
  INVX1 U7508 ( .A(n1558), .Y(n5814) );
  AND2X1 U7509 ( .A(\RF[9][2] ), .B(n10720), .Y(n1546) );
  INVX1 U7510 ( .A(n1546), .Y(n5815) );
  AND2X1 U7511 ( .A(\RF[10][39] ), .B(n10721), .Y(n1518) );
  INVX1 U7512 ( .A(n1518), .Y(n5816) );
  AND2X1 U7513 ( .A(\RF[10][27] ), .B(n10722), .Y(n1506) );
  INVX1 U7514 ( .A(n1506), .Y(n5817) );
  AND2X1 U7515 ( .A(\RF[10][15] ), .B(n10722), .Y(n1494) );
  INVX1 U7516 ( .A(n1494), .Y(n5818) );
  AND2X1 U7517 ( .A(\RF[10][3] ), .B(n10722), .Y(n1482) );
  INVX1 U7518 ( .A(n1482), .Y(n5819) );
  AND2X1 U7519 ( .A(\RF[11][40] ), .B(n10723), .Y(n1454) );
  INVX1 U7520 ( .A(n1454), .Y(n5820) );
  AND2X1 U7521 ( .A(\RF[11][28] ), .B(n10724), .Y(n1442) );
  INVX1 U7522 ( .A(n1442), .Y(n5821) );
  AND2X1 U7523 ( .A(\RF[11][16] ), .B(n10724), .Y(n1430) );
  INVX1 U7524 ( .A(n1430), .Y(n5822) );
  AND2X1 U7525 ( .A(\RF[11][4] ), .B(n10724), .Y(n1418) );
  INVX1 U7526 ( .A(n1418), .Y(n5823) );
  AND2X1 U7527 ( .A(\RF[12][44] ), .B(n10725), .Y(n1393) );
  INVX1 U7528 ( .A(n1393), .Y(n5824) );
  AND2X1 U7529 ( .A(\RF[12][33] ), .B(n10726), .Y(n1382) );
  INVX1 U7530 ( .A(n1382), .Y(n5825) );
  AND2X1 U7531 ( .A(\RF[12][21] ), .B(n10726), .Y(n1370) );
  INVX1 U7532 ( .A(n1370), .Y(n5826) );
  AND2X1 U7533 ( .A(\RF[12][9] ), .B(n10726), .Y(n1358) );
  INVX1 U7534 ( .A(n1358), .Y(n5827) );
  AND2X1 U7535 ( .A(\RF[13][63] ), .B(n10727), .Y(n1347) );
  INVX1 U7536 ( .A(n1347), .Y(n5828) );
  AND2X1 U7537 ( .A(\RF[13][34] ), .B(n10728), .Y(n1318) );
  INVX1 U7538 ( .A(n1318), .Y(n5829) );
  AND2X1 U7539 ( .A(\RF[13][22] ), .B(n10727), .Y(n1306) );
  INVX1 U7540 ( .A(n1306), .Y(n5830) );
  AND2X1 U7541 ( .A(\RF[13][10] ), .B(n10728), .Y(n1294) );
  INVX1 U7542 ( .A(n1294), .Y(n5831) );
  AND2X1 U7543 ( .A(\RF[14][56] ), .B(n10730), .Y(n1275) );
  INVX1 U7544 ( .A(n1275), .Y(n5832) );
  AND2X1 U7545 ( .A(\RF[14][35] ), .B(n10730), .Y(n1254) );
  INVX1 U7546 ( .A(n1254), .Y(n5833) );
  AND2X1 U7547 ( .A(\RF[14][23] ), .B(n10730), .Y(n1242) );
  INVX1 U7548 ( .A(n1242), .Y(n5834) );
  AND2X1 U7549 ( .A(\RF[14][11] ), .B(n10730), .Y(n1230) );
  INVX1 U7550 ( .A(n1230), .Y(n5835) );
  AND2X1 U7551 ( .A(\RF[15][59] ), .B(n10731), .Y(n1212) );
  INVX1 U7552 ( .A(n1212), .Y(n5836) );
  AND2X1 U7553 ( .A(\RF[15][42] ), .B(n10732), .Y(n1195) );
  INVX1 U7554 ( .A(n1195), .Y(n5837) );
  AND2X1 U7555 ( .A(\RF[15][36] ), .B(n10732), .Y(n1189) );
  INVX1 U7556 ( .A(n1189), .Y(n5838) );
  AND2X1 U7557 ( .A(\RF[15][12] ), .B(n10732), .Y(n1165) );
  INVX1 U7558 ( .A(n1165), .Y(n5839) );
  AND2X1 U7559 ( .A(\RF[16][41] ), .B(n10733), .Y(n1129) );
  INVX1 U7560 ( .A(n1129), .Y(n5840) );
  AND2X1 U7561 ( .A(\RF[16][29] ), .B(n10734), .Y(n1117) );
  INVX1 U7562 ( .A(n1117), .Y(n5841) );
  AND2X1 U7563 ( .A(\RF[16][17] ), .B(n10734), .Y(n1105) );
  INVX1 U7564 ( .A(n1105), .Y(n5842) );
  AND2X1 U7565 ( .A(\RF[16][5] ), .B(n10733), .Y(n1093) );
  INVX1 U7566 ( .A(n1093), .Y(n5843) );
  AND2X1 U7567 ( .A(\RF[17][38] ), .B(n10736), .Y(n1061) );
  INVX1 U7568 ( .A(n1061), .Y(n5844) );
  AND2X1 U7569 ( .A(\RF[17][30] ), .B(n10735), .Y(n1053) );
  INVX1 U7570 ( .A(n1053), .Y(n5845) );
  AND2X1 U7571 ( .A(\RF[17][18] ), .B(n10736), .Y(n1041) );
  INVX1 U7572 ( .A(n1041), .Y(n5846) );
  AND2X1 U7573 ( .A(\RF[17][6] ), .B(n10736), .Y(n1029) );
  INVX1 U7574 ( .A(n1029), .Y(n5847) );
  AND2X1 U7575 ( .A(\RF[18][43] ), .B(n10737), .Y(n1001) );
  INVX1 U7576 ( .A(n1001), .Y(n5848) );
  AND2X1 U7577 ( .A(\RF[18][31] ), .B(n10738), .Y(n989) );
  INVX1 U7578 ( .A(n989), .Y(n5849) );
  AND2X1 U7579 ( .A(\RF[18][19] ), .B(n10738), .Y(n977) );
  INVX1 U7580 ( .A(n977), .Y(n5850) );
  AND2X1 U7581 ( .A(\RF[18][7] ), .B(n10738), .Y(n965) );
  INVX1 U7582 ( .A(n965), .Y(n5851) );
  AND2X1 U7583 ( .A(\RF[19][47] ), .B(n10739), .Y(n940) );
  INVX1 U7584 ( .A(n940), .Y(n5852) );
  AND2X1 U7585 ( .A(\RF[19][25] ), .B(n10740), .Y(n918) );
  INVX1 U7586 ( .A(n918), .Y(n5853) );
  AND2X1 U7587 ( .A(\RF[19][20] ), .B(n10740), .Y(n913) );
  INVX1 U7588 ( .A(n913), .Y(n5854) );
  AND2X1 U7589 ( .A(\RF[19][8] ), .B(n10740), .Y(n901) );
  INVX1 U7590 ( .A(n901), .Y(n5855) );
  AND2X1 U7591 ( .A(\RF[20][45] ), .B(n10742), .Y(n873) );
  INVX1 U7592 ( .A(n873), .Y(n5856) );
  AND2X1 U7593 ( .A(\RF[20][32] ), .B(n10741), .Y(n860) );
  INVX1 U7594 ( .A(n860), .Y(n5857) );
  AND2X1 U7595 ( .A(\RF[20][13] ), .B(n10742), .Y(n841) );
  INVX1 U7596 ( .A(n841), .Y(n5858) );
  AND2X1 U7597 ( .A(\RF[20][1] ), .B(n10742), .Y(n829) );
  INVX1 U7598 ( .A(n829), .Y(n5859) );
  AND2X1 U7599 ( .A(\RF[20][0] ), .B(n10741), .Y(n828) );
  INVX1 U7600 ( .A(n828), .Y(n5860) );
  AND2X1 U7601 ( .A(\RF[21][37] ), .B(n10743), .Y(n800) );
  INVX1 U7602 ( .A(n800), .Y(n5861) );
  AND2X1 U7603 ( .A(\RF[21][26] ), .B(n10744), .Y(n789) );
  INVX1 U7604 ( .A(n789), .Y(n5862) );
  AND2X1 U7605 ( .A(\RF[21][14] ), .B(n10744), .Y(n777) );
  INVX1 U7606 ( .A(n777), .Y(n5863) );
  AND2X1 U7607 ( .A(\RF[21][2] ), .B(n10744), .Y(n765) );
  INVX1 U7608 ( .A(n765), .Y(n5864) );
  AND2X1 U7609 ( .A(\RF[22][39] ), .B(n10745), .Y(n737) );
  INVX1 U7610 ( .A(n737), .Y(n5865) );
  AND2X1 U7611 ( .A(\RF[22][27] ), .B(n10746), .Y(n725) );
  INVX1 U7612 ( .A(n725), .Y(n5866) );
  AND2X1 U7613 ( .A(\RF[22][15] ), .B(n10746), .Y(n713) );
  INVX1 U7614 ( .A(n713), .Y(n5867) );
  AND2X1 U7615 ( .A(\RF[22][3] ), .B(n10746), .Y(n701) );
  INVX1 U7616 ( .A(n701), .Y(n5868) );
  AND2X1 U7617 ( .A(\RF[23][40] ), .B(n10747), .Y(n672) );
  INVX1 U7618 ( .A(n672), .Y(n5869) );
  AND2X1 U7619 ( .A(\RF[23][28] ), .B(n10748), .Y(n660) );
  INVX1 U7620 ( .A(n660), .Y(n5870) );
  AND2X1 U7621 ( .A(\RF[23][16] ), .B(n10748), .Y(n648) );
  INVX1 U7622 ( .A(n648), .Y(n5871) );
  AND2X1 U7623 ( .A(\RF[23][4] ), .B(n10748), .Y(n636) );
  INVX1 U7624 ( .A(n636), .Y(n5872) );
  AND2X1 U7625 ( .A(\RF[24][41] ), .B(n10749), .Y(n606) );
  INVX1 U7626 ( .A(n606), .Y(n5873) );
  AND2X1 U7627 ( .A(\RF[24][29] ), .B(n10750), .Y(n594) );
  INVX1 U7628 ( .A(n594), .Y(n5874) );
  AND2X1 U7629 ( .A(\RF[24][17] ), .B(n10750), .Y(n582) );
  INVX1 U7630 ( .A(n582), .Y(n5875) );
  AND2X1 U7631 ( .A(\RF[24][5] ), .B(n10749), .Y(n570) );
  INVX1 U7632 ( .A(n570), .Y(n5876) );
  AND2X1 U7633 ( .A(\RF[25][38] ), .B(n10752), .Y(n537) );
  INVX1 U7634 ( .A(n537), .Y(n5877) );
  AND2X1 U7635 ( .A(\RF[25][30] ), .B(n10751), .Y(n529) );
  INVX1 U7636 ( .A(n529), .Y(n5878) );
  AND2X1 U7637 ( .A(\RF[25][18] ), .B(n10752), .Y(n517) );
  INVX1 U7638 ( .A(n517), .Y(n5879) );
  AND2X1 U7639 ( .A(\RF[25][6] ), .B(n10752), .Y(n505) );
  INVX1 U7640 ( .A(n505), .Y(n5880) );
  AND2X1 U7641 ( .A(\RF[26][43] ), .B(n10753), .Y(n476) );
  INVX1 U7642 ( .A(n476), .Y(n5881) );
  AND2X1 U7643 ( .A(\RF[26][31] ), .B(n10754), .Y(n464) );
  INVX1 U7644 ( .A(n464), .Y(n5882) );
  AND2X1 U7645 ( .A(\RF[26][19] ), .B(n10754), .Y(n452) );
  INVX1 U7646 ( .A(n452), .Y(n5883) );
  AND2X1 U7647 ( .A(\RF[26][7] ), .B(n10754), .Y(n440) );
  INVX1 U7648 ( .A(n440), .Y(n5884) );
  AND2X1 U7649 ( .A(\RF[27][47] ), .B(n10755), .Y(n414) );
  INVX1 U7650 ( .A(n414), .Y(n5885) );
  AND2X1 U7651 ( .A(\RF[27][25] ), .B(n10756), .Y(n392) );
  INVX1 U7652 ( .A(n392), .Y(n5886) );
  AND2X1 U7653 ( .A(\RF[27][20] ), .B(n10756), .Y(n387) );
  INVX1 U7654 ( .A(n387), .Y(n5887) );
  AND2X1 U7655 ( .A(\RF[27][8] ), .B(n10756), .Y(n375) );
  INVX1 U7656 ( .A(n375), .Y(n5888) );
  AND2X1 U7657 ( .A(\RF[28][45] ), .B(n10758), .Y(n346) );
  INVX1 U7658 ( .A(n346), .Y(n5889) );
  AND2X1 U7659 ( .A(\RF[28][32] ), .B(n10757), .Y(n333) );
  INVX1 U7660 ( .A(n333), .Y(n5890) );
  AND2X1 U7661 ( .A(\RF[28][13] ), .B(n10758), .Y(n314) );
  INVX1 U7662 ( .A(n314), .Y(n5891) );
  AND2X1 U7663 ( .A(\RF[28][1] ), .B(n10758), .Y(n302) );
  INVX1 U7664 ( .A(n302), .Y(n5892) );
  AND2X1 U7665 ( .A(\RF[28][0] ), .B(n10757), .Y(n301) );
  INVX1 U7666 ( .A(n301), .Y(n5893) );
  AND2X1 U7667 ( .A(\RF[29][37] ), .B(n10759), .Y(n272) );
  INVX1 U7668 ( .A(n272), .Y(n5894) );
  AND2X1 U7669 ( .A(\RF[29][26] ), .B(n10760), .Y(n261) );
  INVX1 U7670 ( .A(n261), .Y(n5895) );
  AND2X1 U7671 ( .A(\RF[29][14] ), .B(n10760), .Y(n249) );
  INVX1 U7672 ( .A(n249), .Y(n5896) );
  AND2X1 U7673 ( .A(\RF[29][2] ), .B(n10760), .Y(n237) );
  INVX1 U7674 ( .A(n237), .Y(n5897) );
  AND2X1 U7675 ( .A(\RF[30][39] ), .B(n10761), .Y(n208) );
  INVX1 U7676 ( .A(n208), .Y(n5898) );
  AND2X1 U7677 ( .A(\RF[30][27] ), .B(n10762), .Y(n196) );
  INVX1 U7678 ( .A(n196), .Y(n5899) );
  AND2X1 U7679 ( .A(\RF[30][15] ), .B(n10762), .Y(n184) );
  INVX1 U7680 ( .A(n184), .Y(n5900) );
  AND2X1 U7681 ( .A(\RF[30][3] ), .B(n10762), .Y(n172) );
  INVX1 U7682 ( .A(n172), .Y(n5901) );
  AND2X1 U7683 ( .A(\RF[31][40] ), .B(n10763), .Y(n119) );
  INVX1 U7684 ( .A(n119), .Y(n5902) );
  AND2X1 U7685 ( .A(\RF[31][28] ), .B(n10764), .Y(n95) );
  INVX1 U7686 ( .A(n95), .Y(n5903) );
  AND2X1 U7687 ( .A(\RF[31][16] ), .B(n10764), .Y(n71) );
  INVX1 U7688 ( .A(n71), .Y(n5904) );
  AND2X1 U7689 ( .A(\RF[31][4] ), .B(n10764), .Y(n47) );
  INVX1 U7690 ( .A(n47), .Y(n5905) );
  BUFX2 U7691 ( .A(n167), .Y(n5906) );
  AND2X1 U7692 ( .A(\RF[0][63] ), .B(n10701), .Y(n2193) );
  INVX1 U7693 ( .A(n2193), .Y(n5907) );
  AND2X1 U7694 ( .A(\RF[0][34] ), .B(n10702), .Y(n2164) );
  INVX1 U7695 ( .A(n2164), .Y(n5908) );
  AND2X1 U7696 ( .A(\RF[0][22] ), .B(n10702), .Y(n2152) );
  INVX1 U7697 ( .A(n2152), .Y(n5909) );
  AND2X1 U7698 ( .A(\RF[0][10] ), .B(n10702), .Y(n2140) );
  INVX1 U7699 ( .A(n2140), .Y(n5910) );
  AND2X1 U7700 ( .A(\RF[1][44] ), .B(n10704), .Y(n2109) );
  INVX1 U7701 ( .A(n2109), .Y(n5911) );
  AND2X1 U7702 ( .A(\RF[1][33] ), .B(n10704), .Y(n2098) );
  INVX1 U7703 ( .A(n2098), .Y(n5912) );
  AND2X1 U7704 ( .A(\RF[1][21] ), .B(n10704), .Y(n2086) );
  INVX1 U7705 ( .A(n2086), .Y(n5913) );
  AND2X1 U7706 ( .A(\RF[1][9] ), .B(n10704), .Y(n2074) );
  INVX1 U7707 ( .A(n2074), .Y(n5914) );
  AND2X1 U7708 ( .A(\RF[2][59] ), .B(n10705), .Y(n2059) );
  INVX1 U7709 ( .A(n2059), .Y(n5915) );
  AND2X1 U7710 ( .A(\RF[2][42] ), .B(n10706), .Y(n2042) );
  INVX1 U7711 ( .A(n2042), .Y(n5916) );
  AND2X1 U7712 ( .A(\RF[2][36] ), .B(n10705), .Y(n2036) );
  INVX1 U7713 ( .A(n2036), .Y(n5917) );
  AND2X1 U7714 ( .A(\RF[2][12] ), .B(n10706), .Y(n2012) );
  INVX1 U7715 ( .A(n2012), .Y(n5918) );
  AND2X1 U7716 ( .A(\RF[3][56] ), .B(n10708), .Y(n1991) );
  INVX1 U7717 ( .A(n1991), .Y(n5919) );
  AND2X1 U7718 ( .A(\RF[3][35] ), .B(n10707), .Y(n1970) );
  INVX1 U7719 ( .A(n1970), .Y(n5920) );
  AND2X1 U7720 ( .A(\RF[3][23] ), .B(n10708), .Y(n1958) );
  INVX1 U7721 ( .A(n1958), .Y(n5921) );
  AND2X1 U7722 ( .A(\RF[3][11] ), .B(n10708), .Y(n1946) );
  INVX1 U7723 ( .A(n1946), .Y(n5922) );
  AND2X1 U7724 ( .A(\RF[4][38] ), .B(n10710), .Y(n1908) );
  INVX1 U7725 ( .A(n1908), .Y(n5923) );
  AND2X1 U7726 ( .A(\RF[4][30] ), .B(n10710), .Y(n1900) );
  INVX1 U7727 ( .A(n1900), .Y(n5924) );
  AND2X1 U7728 ( .A(\RF[4][18] ), .B(n10710), .Y(n1888) );
  INVX1 U7729 ( .A(n1888), .Y(n5925) );
  AND2X1 U7730 ( .A(\RF[4][6] ), .B(n10710), .Y(n1876) );
  INVX1 U7731 ( .A(n1876), .Y(n5926) );
  AND2X1 U7732 ( .A(\RF[5][41] ), .B(n10712), .Y(n1846) );
  INVX1 U7733 ( .A(n1846), .Y(n5927) );
  AND2X1 U7734 ( .A(\RF[5][29] ), .B(n10712), .Y(n1834) );
  INVX1 U7735 ( .A(n1834), .Y(n5928) );
  AND2X1 U7736 ( .A(\RF[5][17] ), .B(n10712), .Y(n1822) );
  INVX1 U7737 ( .A(n1822), .Y(n5929) );
  AND2X1 U7738 ( .A(\RF[5][5] ), .B(n10711), .Y(n1810) );
  INVX1 U7739 ( .A(n1810), .Y(n5930) );
  AND2X1 U7740 ( .A(\RF[6][47] ), .B(n10714), .Y(n1787) );
  INVX1 U7741 ( .A(n1787), .Y(n5931) );
  AND2X1 U7742 ( .A(\RF[6][25] ), .B(n10714), .Y(n1765) );
  INVX1 U7743 ( .A(n1765), .Y(n5932) );
  AND2X1 U7744 ( .A(\RF[6][20] ), .B(n10714), .Y(n1760) );
  INVX1 U7745 ( .A(n1760), .Y(n5933) );
  AND2X1 U7746 ( .A(\RF[6][8] ), .B(n10713), .Y(n1748) );
  INVX1 U7747 ( .A(n1748), .Y(n5934) );
  AND2X1 U7748 ( .A(\RF[7][43] ), .B(n10716), .Y(n1717) );
  INVX1 U7749 ( .A(n1717), .Y(n5935) );
  AND2X1 U7750 ( .A(\RF[7][31] ), .B(n10716), .Y(n1705) );
  INVX1 U7751 ( .A(n1705), .Y(n5936) );
  AND2X1 U7752 ( .A(\RF[7][19] ), .B(n10716), .Y(n1693) );
  INVX1 U7753 ( .A(n1693), .Y(n5937) );
  AND2X1 U7754 ( .A(\RF[7][7] ), .B(n10715), .Y(n1681) );
  INVX1 U7755 ( .A(n1681), .Y(n5938) );
  AND2X1 U7756 ( .A(\RF[8][37] ), .B(n10718), .Y(n1646) );
  INVX1 U7757 ( .A(n1646), .Y(n5939) );
  AND2X1 U7758 ( .A(\RF[8][26] ), .B(n10718), .Y(n1635) );
  INVX1 U7759 ( .A(n1635), .Y(n5940) );
  AND2X1 U7760 ( .A(\RF[8][14] ), .B(n10718), .Y(n1623) );
  INVX1 U7761 ( .A(n1623), .Y(n5941) );
  AND2X1 U7762 ( .A(\RF[8][2] ), .B(n10717), .Y(n1611) );
  INVX1 U7763 ( .A(n1611), .Y(n5942) );
  AND2X1 U7764 ( .A(\RF[9][45] ), .B(n10720), .Y(n1589) );
  INVX1 U7765 ( .A(n1589), .Y(n5943) );
  AND2X1 U7766 ( .A(\RF[9][32] ), .B(n10720), .Y(n1576) );
  INVX1 U7767 ( .A(n1576), .Y(n5944) );
  AND2X1 U7768 ( .A(\RF[9][13] ), .B(n10720), .Y(n1557) );
  INVX1 U7769 ( .A(n1557), .Y(n5945) );
  AND2X1 U7770 ( .A(\RF[9][1] ), .B(n10719), .Y(n1545) );
  INVX1 U7771 ( .A(n1545), .Y(n5946) );
  AND2X1 U7772 ( .A(\RF[9][0] ), .B(n10719), .Y(n1544) );
  INVX1 U7773 ( .A(n1544), .Y(n5947) );
  AND2X1 U7774 ( .A(\RF[10][40] ), .B(n10722), .Y(n1519) );
  INVX1 U7775 ( .A(n1519), .Y(n5948) );
  AND2X1 U7776 ( .A(\RF[10][28] ), .B(n10722), .Y(n1507) );
  INVX1 U7777 ( .A(n1507), .Y(n5949) );
  AND2X1 U7778 ( .A(\RF[10][16] ), .B(n10722), .Y(n1495) );
  INVX1 U7779 ( .A(n1495), .Y(n5950) );
  AND2X1 U7780 ( .A(\RF[10][4] ), .B(n10721), .Y(n1483) );
  INVX1 U7781 ( .A(n1483), .Y(n5951) );
  AND2X1 U7782 ( .A(\RF[11][39] ), .B(n10724), .Y(n1453) );
  INVX1 U7783 ( .A(n1453), .Y(n5952) );
  AND2X1 U7784 ( .A(\RF[11][27] ), .B(n10724), .Y(n1441) );
  INVX1 U7785 ( .A(n1441), .Y(n5953) );
  AND2X1 U7786 ( .A(\RF[11][15] ), .B(n10724), .Y(n1429) );
  INVX1 U7787 ( .A(n1429), .Y(n5954) );
  AND2X1 U7788 ( .A(\RF[11][3] ), .B(n10723), .Y(n1417) );
  INVX1 U7789 ( .A(n1417), .Y(n5955) );
  AND2X1 U7790 ( .A(\RF[12][63] ), .B(n10725), .Y(n1412) );
  INVX1 U7791 ( .A(n1412), .Y(n5956) );
  AND2X1 U7792 ( .A(\RF[12][34] ), .B(n10726), .Y(n1383) );
  INVX1 U7793 ( .A(n1383), .Y(n5957) );
  AND2X1 U7794 ( .A(\RF[12][22] ), .B(n10726), .Y(n1371) );
  INVX1 U7795 ( .A(n1371), .Y(n5958) );
  AND2X1 U7796 ( .A(\RF[12][10] ), .B(n10726), .Y(n1359) );
  INVX1 U7797 ( .A(n1359), .Y(n5959) );
  AND2X1 U7798 ( .A(\RF[13][44] ), .B(n10728), .Y(n1328) );
  INVX1 U7799 ( .A(n1328), .Y(n5960) );
  AND2X1 U7800 ( .A(\RF[13][33] ), .B(n10728), .Y(n1317) );
  INVX1 U7801 ( .A(n1317), .Y(n5961) );
  AND2X1 U7802 ( .A(\RF[13][21] ), .B(n10728), .Y(n1305) );
  INVX1 U7803 ( .A(n1305), .Y(n5962) );
  AND2X1 U7804 ( .A(\RF[13][9] ), .B(n10728), .Y(n1293) );
  INVX1 U7805 ( .A(n1293), .Y(n5963) );
  AND2X1 U7806 ( .A(\RF[14][59] ), .B(n10729), .Y(n1278) );
  INVX1 U7807 ( .A(n1278), .Y(n5964) );
  AND2X1 U7808 ( .A(\RF[14][42] ), .B(n10730), .Y(n1261) );
  INVX1 U7809 ( .A(n1261), .Y(n5965) );
  AND2X1 U7810 ( .A(\RF[14][36] ), .B(n10729), .Y(n1255) );
  INVX1 U7811 ( .A(n1255), .Y(n5966) );
  AND2X1 U7812 ( .A(\RF[14][12] ), .B(n10730), .Y(n1231) );
  INVX1 U7813 ( .A(n1231), .Y(n5967) );
  AND2X1 U7814 ( .A(\RF[15][56] ), .B(n10732), .Y(n1209) );
  INVX1 U7815 ( .A(n1209), .Y(n5968) );
  AND2X1 U7816 ( .A(\RF[15][35] ), .B(n10731), .Y(n1188) );
  INVX1 U7817 ( .A(n1188), .Y(n5969) );
  AND2X1 U7818 ( .A(\RF[15][23] ), .B(n10732), .Y(n1176) );
  INVX1 U7819 ( .A(n1176), .Y(n5970) );
  AND2X1 U7820 ( .A(\RF[15][11] ), .B(n10732), .Y(n1164) );
  INVX1 U7821 ( .A(n1164), .Y(n5971) );
  AND2X1 U7822 ( .A(\RF[16][38] ), .B(n10734), .Y(n1126) );
  INVX1 U7823 ( .A(n1126), .Y(n5972) );
  AND2X1 U7824 ( .A(\RF[16][30] ), .B(n10734), .Y(n1118) );
  INVX1 U7825 ( .A(n1118), .Y(n5973) );
  AND2X1 U7826 ( .A(\RF[16][18] ), .B(n10734), .Y(n1106) );
  INVX1 U7827 ( .A(n1106), .Y(n5974) );
  AND2X1 U7828 ( .A(\RF[16][6] ), .B(n10734), .Y(n1094) );
  INVX1 U7829 ( .A(n1094), .Y(n5975) );
  AND2X1 U7830 ( .A(\RF[17][41] ), .B(n10736), .Y(n1064) );
  INVX1 U7831 ( .A(n1064), .Y(n5976) );
  AND2X1 U7832 ( .A(\RF[17][29] ), .B(n10736), .Y(n1052) );
  INVX1 U7833 ( .A(n1052), .Y(n5977) );
  AND2X1 U7834 ( .A(\RF[17][17] ), .B(n10736), .Y(n1040) );
  INVX1 U7835 ( .A(n1040), .Y(n5978) );
  AND2X1 U7836 ( .A(\RF[17][5] ), .B(n10735), .Y(n1028) );
  INVX1 U7837 ( .A(n1028), .Y(n5979) );
  AND2X1 U7838 ( .A(\RF[18][47] ), .B(n10738), .Y(n1005) );
  INVX1 U7839 ( .A(n1005), .Y(n5980) );
  AND2X1 U7840 ( .A(\RF[18][25] ), .B(n10738), .Y(n983) );
  INVX1 U7841 ( .A(n983), .Y(n5981) );
  AND2X1 U7842 ( .A(\RF[18][20] ), .B(n10738), .Y(n978) );
  INVX1 U7843 ( .A(n978), .Y(n5982) );
  AND2X1 U7844 ( .A(\RF[18][8] ), .B(n10737), .Y(n966) );
  INVX1 U7845 ( .A(n966), .Y(n5983) );
  AND2X1 U7846 ( .A(\RF[19][43] ), .B(n10740), .Y(n936) );
  INVX1 U7847 ( .A(n936), .Y(n5984) );
  AND2X1 U7848 ( .A(\RF[19][31] ), .B(n10740), .Y(n924) );
  INVX1 U7849 ( .A(n924), .Y(n5985) );
  AND2X1 U7850 ( .A(\RF[19][19] ), .B(n10740), .Y(n912) );
  INVX1 U7851 ( .A(n912), .Y(n5986) );
  AND2X1 U7852 ( .A(\RF[19][7] ), .B(n10739), .Y(n900) );
  INVX1 U7853 ( .A(n900), .Y(n5987) );
  AND2X1 U7854 ( .A(\RF[20][37] ), .B(n10742), .Y(n865) );
  INVX1 U7855 ( .A(n865), .Y(n5988) );
  AND2X1 U7856 ( .A(\RF[20][26] ), .B(n10742), .Y(n854) );
  INVX1 U7857 ( .A(n854), .Y(n5989) );
  AND2X1 U7858 ( .A(\RF[20][14] ), .B(n10742), .Y(n842) );
  INVX1 U7859 ( .A(n842), .Y(n5990) );
  AND2X1 U7860 ( .A(\RF[20][2] ), .B(n10741), .Y(n830) );
  INVX1 U7861 ( .A(n830), .Y(n5991) );
  AND2X1 U7862 ( .A(\RF[21][45] ), .B(n10744), .Y(n808) );
  INVX1 U7863 ( .A(n808), .Y(n5992) );
  AND2X1 U7864 ( .A(\RF[21][32] ), .B(n10744), .Y(n795) );
  INVX1 U7865 ( .A(n795), .Y(n5993) );
  AND2X1 U7866 ( .A(\RF[21][13] ), .B(n10744), .Y(n776) );
  INVX1 U7867 ( .A(n776), .Y(n5994) );
  AND2X1 U7868 ( .A(\RF[21][1] ), .B(n10743), .Y(n764) );
  INVX1 U7869 ( .A(n764), .Y(n5995) );
  AND2X1 U7870 ( .A(\RF[21][0] ), .B(n10743), .Y(n763) );
  INVX1 U7871 ( .A(n763), .Y(n5996) );
  AND2X1 U7872 ( .A(\RF[22][40] ), .B(n10746), .Y(n738) );
  INVX1 U7873 ( .A(n738), .Y(n5997) );
  AND2X1 U7874 ( .A(\RF[22][28] ), .B(n10746), .Y(n726) );
  INVX1 U7875 ( .A(n726), .Y(n5998) );
  AND2X1 U7876 ( .A(\RF[22][16] ), .B(n10746), .Y(n714) );
  INVX1 U7877 ( .A(n714), .Y(n5999) );
  AND2X1 U7878 ( .A(\RF[22][4] ), .B(n10745), .Y(n702) );
  INVX1 U7879 ( .A(n702), .Y(n6000) );
  AND2X1 U7880 ( .A(\RF[23][39] ), .B(n10748), .Y(n671) );
  INVX1 U7881 ( .A(n671), .Y(n6001) );
  AND2X1 U7882 ( .A(\RF[23][27] ), .B(n10748), .Y(n659) );
  INVX1 U7883 ( .A(n659), .Y(n6002) );
  AND2X1 U7884 ( .A(\RF[23][15] ), .B(n10748), .Y(n647) );
  INVX1 U7885 ( .A(n647), .Y(n6003) );
  AND2X1 U7886 ( .A(\RF[23][3] ), .B(n10747), .Y(n635) );
  INVX1 U7887 ( .A(n635), .Y(n6004) );
  AND2X1 U7888 ( .A(\RF[24][38] ), .B(n10750), .Y(n603) );
  INVX1 U7889 ( .A(n603), .Y(n6005) );
  AND2X1 U7890 ( .A(\RF[24][30] ), .B(n10750), .Y(n595) );
  INVX1 U7891 ( .A(n595), .Y(n6006) );
  AND2X1 U7892 ( .A(\RF[24][18] ), .B(n10750), .Y(n583) );
  INVX1 U7893 ( .A(n583), .Y(n6007) );
  AND2X1 U7894 ( .A(\RF[24][6] ), .B(n10750), .Y(n571) );
  INVX1 U7895 ( .A(n571), .Y(n6008) );
  AND2X1 U7896 ( .A(\RF[25][41] ), .B(n10752), .Y(n540) );
  INVX1 U7897 ( .A(n540), .Y(n6009) );
  AND2X1 U7898 ( .A(\RF[25][29] ), .B(n10752), .Y(n528) );
  INVX1 U7899 ( .A(n528), .Y(n6010) );
  AND2X1 U7900 ( .A(\RF[25][17] ), .B(n10752), .Y(n516) );
  INVX1 U7901 ( .A(n516), .Y(n6011) );
  AND2X1 U7902 ( .A(\RF[25][5] ), .B(n10751), .Y(n504) );
  INVX1 U7903 ( .A(n504), .Y(n6012) );
  AND2X1 U7904 ( .A(\RF[26][47] ), .B(n10754), .Y(n480) );
  INVX1 U7905 ( .A(n480), .Y(n6013) );
  AND2X1 U7906 ( .A(\RF[26][25] ), .B(n10754), .Y(n458) );
  INVX1 U7907 ( .A(n458), .Y(n6014) );
  AND2X1 U7908 ( .A(\RF[26][20] ), .B(n10754), .Y(n453) );
  INVX1 U7909 ( .A(n453), .Y(n6015) );
  AND2X1 U7910 ( .A(\RF[26][8] ), .B(n10753), .Y(n441) );
  INVX1 U7911 ( .A(n441), .Y(n6016) );
  AND2X1 U7912 ( .A(\RF[27][43] ), .B(n10756), .Y(n410) );
  INVX1 U7913 ( .A(n410), .Y(n6017) );
  AND2X1 U7914 ( .A(\RF[27][31] ), .B(n10756), .Y(n398) );
  INVX1 U7915 ( .A(n398), .Y(n6018) );
  AND2X1 U7916 ( .A(\RF[27][19] ), .B(n10756), .Y(n386) );
  INVX1 U7917 ( .A(n386), .Y(n6019) );
  AND2X1 U7918 ( .A(\RF[27][7] ), .B(n10755), .Y(n374) );
  INVX1 U7919 ( .A(n374), .Y(n6020) );
  AND2X1 U7920 ( .A(\RF[28][37] ), .B(n10758), .Y(n338) );
  INVX1 U7921 ( .A(n338), .Y(n6021) );
  AND2X1 U7922 ( .A(\RF[28][26] ), .B(n10758), .Y(n327) );
  INVX1 U7923 ( .A(n327), .Y(n6022) );
  AND2X1 U7924 ( .A(\RF[28][14] ), .B(n10758), .Y(n315) );
  INVX1 U7925 ( .A(n315), .Y(n6023) );
  AND2X1 U7926 ( .A(\RF[28][2] ), .B(n10757), .Y(n303) );
  INVX1 U7927 ( .A(n303), .Y(n6024) );
  AND2X1 U7928 ( .A(\RF[29][45] ), .B(n10760), .Y(n280) );
  INVX1 U7929 ( .A(n280), .Y(n6025) );
  AND2X1 U7930 ( .A(\RF[29][32] ), .B(n10760), .Y(n267) );
  INVX1 U7931 ( .A(n267), .Y(n6026) );
  AND2X1 U7932 ( .A(\RF[29][13] ), .B(n10760), .Y(n248) );
  INVX1 U7933 ( .A(n248), .Y(n6027) );
  AND2X1 U7934 ( .A(\RF[29][1] ), .B(n10759), .Y(n236) );
  INVX1 U7935 ( .A(n236), .Y(n6028) );
  AND2X1 U7936 ( .A(\RF[29][0] ), .B(n10759), .Y(n235) );
  INVX1 U7937 ( .A(n235), .Y(n6029) );
  AND2X1 U7938 ( .A(\RF[30][40] ), .B(n10762), .Y(n209) );
  INVX1 U7939 ( .A(n209), .Y(n6030) );
  AND2X1 U7940 ( .A(\RF[30][28] ), .B(n10762), .Y(n197) );
  INVX1 U7941 ( .A(n197), .Y(n6031) );
  AND2X1 U7942 ( .A(\RF[30][16] ), .B(n10762), .Y(n185) );
  INVX1 U7943 ( .A(n185), .Y(n6032) );
  AND2X1 U7944 ( .A(\RF[30][4] ), .B(n10761), .Y(n173) );
  INVX1 U7945 ( .A(n173), .Y(n6033) );
  AND2X1 U7946 ( .A(\RF[31][39] ), .B(n10764), .Y(n117) );
  INVX1 U7947 ( .A(n117), .Y(n6034) );
  AND2X1 U7948 ( .A(\RF[31][27] ), .B(n10764), .Y(n93) );
  INVX1 U7949 ( .A(n93), .Y(n6035) );
  AND2X1 U7950 ( .A(\RF[31][15] ), .B(n10764), .Y(n69) );
  INVX1 U7951 ( .A(n69), .Y(n6036) );
  AND2X1 U7952 ( .A(\RF[31][3] ), .B(n10763), .Y(n45) );
  INVX1 U7953 ( .A(n45), .Y(n6037) );
  BUFX2 U7954 ( .A(n1739), .Y(n6038) );
  AND2X1 U7955 ( .A(\RF[0][56] ), .B(n10702), .Y(n2186) );
  INVX1 U7956 ( .A(n2186), .Y(n6039) );
  AND2X1 U7957 ( .A(\RF[0][35] ), .B(n10701), .Y(n2165) );
  INVX1 U7958 ( .A(n2165), .Y(n6040) );
  AND2X1 U7959 ( .A(\RF[0][23] ), .B(n10701), .Y(n2153) );
  INVX1 U7960 ( .A(n2153), .Y(n6041) );
  AND2X1 U7961 ( .A(\RF[0][11] ), .B(n10701), .Y(n2141) );
  INVX1 U7962 ( .A(n2141), .Y(n6042) );
  AND2X1 U7963 ( .A(\RF[1][59] ), .B(n10704), .Y(n2124) );
  INVX1 U7964 ( .A(n2124), .Y(n6043) );
  AND2X1 U7965 ( .A(\RF[1][42] ), .B(n10703), .Y(n2107) );
  INVX1 U7966 ( .A(n2107), .Y(n6044) );
  AND2X1 U7967 ( .A(\RF[1][36] ), .B(n10703), .Y(n2101) );
  INVX1 U7968 ( .A(n2101), .Y(n6045) );
  AND2X1 U7969 ( .A(\RF[1][12] ), .B(n10703), .Y(n2077) );
  INVX1 U7970 ( .A(n2077), .Y(n6046) );
  AND2X1 U7971 ( .A(\RF[2][44] ), .B(n10705), .Y(n2044) );
  INVX1 U7972 ( .A(n2044), .Y(n6047) );
  AND2X1 U7973 ( .A(\RF[2][33] ), .B(n10706), .Y(n2033) );
  INVX1 U7974 ( .A(n2033), .Y(n6048) );
  AND2X1 U7975 ( .A(\RF[2][21] ), .B(n10706), .Y(n2021) );
  INVX1 U7976 ( .A(n2021), .Y(n6049) );
  AND2X1 U7977 ( .A(\RF[2][9] ), .B(n10705), .Y(n2009) );
  INVX1 U7978 ( .A(n2009), .Y(n6050) );
  AND2X1 U7979 ( .A(\RF[3][63] ), .B(n10707), .Y(n1998) );
  INVX1 U7980 ( .A(n1998), .Y(n6051) );
  AND2X1 U7981 ( .A(\RF[3][34] ), .B(n10707), .Y(n1969) );
  INVX1 U7982 ( .A(n1969), .Y(n6052) );
  AND2X1 U7983 ( .A(\RF[3][22] ), .B(n10708), .Y(n1957) );
  INVX1 U7984 ( .A(n1957), .Y(n6053) );
  AND2X1 U7985 ( .A(\RF[3][10] ), .B(n10707), .Y(n1945) );
  INVX1 U7986 ( .A(n1945), .Y(n6054) );
  AND2X1 U7987 ( .A(\RF[4][43] ), .B(n10709), .Y(n1913) );
  INVX1 U7988 ( .A(n1913), .Y(n6055) );
  AND2X1 U7989 ( .A(\RF[4][31] ), .B(n10709), .Y(n1901) );
  INVX1 U7990 ( .A(n1901), .Y(n6056) );
  AND2X1 U7991 ( .A(\RF[4][19] ), .B(n10710), .Y(n1889) );
  INVX1 U7992 ( .A(n1889), .Y(n6057) );
  AND2X1 U7993 ( .A(\RF[4][7] ), .B(n10709), .Y(n1877) );
  INVX1 U7994 ( .A(n1877), .Y(n6058) );
  AND2X1 U7995 ( .A(\RF[5][47] ), .B(n10711), .Y(n1852) );
  INVX1 U7996 ( .A(n1852), .Y(n6059) );
  AND2X1 U7997 ( .A(\RF[5][25] ), .B(n10711), .Y(n1830) );
  INVX1 U7998 ( .A(n1830), .Y(n6060) );
  AND2X1 U7999 ( .A(\RF[5][20] ), .B(n10712), .Y(n1825) );
  INVX1 U8000 ( .A(n1825), .Y(n6061) );
  AND2X1 U8001 ( .A(\RF[5][8] ), .B(n10711), .Y(n1813) );
  INVX1 U8002 ( .A(n1813), .Y(n6062) );
  AND2X1 U8003 ( .A(\RF[6][41] ), .B(n10713), .Y(n1781) );
  INVX1 U8004 ( .A(n1781), .Y(n6063) );
  AND2X1 U8005 ( .A(\RF[6][29] ), .B(n10714), .Y(n1769) );
  INVX1 U8006 ( .A(n1769), .Y(n6064) );
  AND2X1 U8007 ( .A(\RF[6][17] ), .B(n10713), .Y(n1757) );
  INVX1 U8008 ( .A(n1757), .Y(n6065) );
  AND2X1 U8009 ( .A(\RF[6][5] ), .B(n10713), .Y(n1745) );
  INVX1 U8010 ( .A(n1745), .Y(n6066) );
  AND2X1 U8011 ( .A(\RF[7][38] ), .B(n10716), .Y(n1712) );
  INVX1 U8012 ( .A(n1712), .Y(n6067) );
  AND2X1 U8013 ( .A(\RF[7][30] ), .B(n10715), .Y(n1704) );
  INVX1 U8014 ( .A(n1704), .Y(n6068) );
  AND2X1 U8015 ( .A(\RF[7][18] ), .B(n10715), .Y(n1692) );
  INVX1 U8016 ( .A(n1692), .Y(n6069) );
  AND2X1 U8017 ( .A(\RF[7][6] ), .B(n10715), .Y(n1680) );
  INVX1 U8018 ( .A(n1680), .Y(n6070) );
  AND2X1 U8019 ( .A(\RF[8][39] ), .B(n10717), .Y(n1648) );
  INVX1 U8020 ( .A(n1648), .Y(n6071) );
  AND2X1 U8021 ( .A(\RF[8][27] ), .B(n10718), .Y(n1636) );
  INVX1 U8022 ( .A(n1636), .Y(n6072) );
  AND2X1 U8023 ( .A(\RF[8][15] ), .B(n10717), .Y(n1624) );
  INVX1 U8024 ( .A(n1624), .Y(n6073) );
  AND2X1 U8025 ( .A(\RF[8][3] ), .B(n10717), .Y(n1612) );
  INVX1 U8026 ( .A(n1612), .Y(n6074) );
  AND2X1 U8027 ( .A(\RF[9][40] ), .B(n10719), .Y(n1584) );
  INVX1 U8028 ( .A(n1584), .Y(n6075) );
  AND2X1 U8029 ( .A(\RF[9][28] ), .B(n10720), .Y(n1572) );
  INVX1 U8030 ( .A(n1572), .Y(n6076) );
  AND2X1 U8031 ( .A(\RF[9][16] ), .B(n10719), .Y(n1560) );
  INVX1 U8032 ( .A(n1560), .Y(n6077) );
  AND2X1 U8033 ( .A(\RF[9][4] ), .B(n10719), .Y(n1548) );
  INVX1 U8034 ( .A(n1548), .Y(n6078) );
  AND2X1 U8035 ( .A(\RF[10][45] ), .B(n10722), .Y(n1524) );
  INVX1 U8036 ( .A(n1524), .Y(n6079) );
  AND2X1 U8037 ( .A(\RF[10][32] ), .B(n10721), .Y(n1511) );
  INVX1 U8038 ( .A(n1511), .Y(n6080) );
  AND2X1 U8039 ( .A(\RF[10][13] ), .B(n10721), .Y(n1492) );
  INVX1 U8040 ( .A(n1492), .Y(n6081) );
  AND2X1 U8041 ( .A(\RF[10][1] ), .B(n10721), .Y(n1480) );
  INVX1 U8042 ( .A(n1480), .Y(n6082) );
  AND2X1 U8043 ( .A(\RF[10][0] ), .B(n10721), .Y(n1479) );
  INVX1 U8044 ( .A(n1479), .Y(n6083) );
  AND2X1 U8045 ( .A(\RF[11][37] ), .B(n10723), .Y(n1451) );
  INVX1 U8046 ( .A(n1451), .Y(n6084) );
  AND2X1 U8047 ( .A(\RF[11][26] ), .B(n10724), .Y(n1440) );
  INVX1 U8048 ( .A(n1440), .Y(n6085) );
  AND2X1 U8049 ( .A(\RF[11][14] ), .B(n10723), .Y(n1428) );
  INVX1 U8050 ( .A(n1428), .Y(n6086) );
  AND2X1 U8051 ( .A(\RF[11][2] ), .B(n10723), .Y(n1416) );
  INVX1 U8052 ( .A(n1416), .Y(n6087) );
  AND2X1 U8053 ( .A(\RF[12][56] ), .B(n10726), .Y(n1405) );
  INVX1 U8054 ( .A(n1405), .Y(n6088) );
  AND2X1 U8055 ( .A(\RF[12][35] ), .B(n10725), .Y(n1384) );
  INVX1 U8056 ( .A(n1384), .Y(n6089) );
  AND2X1 U8057 ( .A(\RF[12][23] ), .B(n10725), .Y(n1372) );
  INVX1 U8058 ( .A(n1372), .Y(n6090) );
  AND2X1 U8059 ( .A(\RF[12][11] ), .B(n10725), .Y(n1360) );
  INVX1 U8060 ( .A(n1360), .Y(n6091) );
  AND2X1 U8061 ( .A(\RF[13][59] ), .B(n10728), .Y(n1343) );
  INVX1 U8062 ( .A(n1343), .Y(n6092) );
  AND2X1 U8063 ( .A(\RF[13][42] ), .B(n10727), .Y(n1326) );
  INVX1 U8064 ( .A(n1326), .Y(n6093) );
  AND2X1 U8065 ( .A(\RF[13][36] ), .B(n10727), .Y(n1320) );
  INVX1 U8066 ( .A(n1320), .Y(n6094) );
  AND2X1 U8067 ( .A(\RF[13][12] ), .B(n10727), .Y(n1296) );
  INVX1 U8068 ( .A(n1296), .Y(n6095) );
  AND2X1 U8069 ( .A(\RF[14][44] ), .B(n10729), .Y(n1263) );
  INVX1 U8070 ( .A(n1263), .Y(n6096) );
  AND2X1 U8071 ( .A(\RF[14][33] ), .B(n10730), .Y(n1252) );
  INVX1 U8072 ( .A(n1252), .Y(n6097) );
  AND2X1 U8073 ( .A(\RF[14][21] ), .B(n10730), .Y(n1240) );
  INVX1 U8074 ( .A(n1240), .Y(n6098) );
  AND2X1 U8075 ( .A(\RF[14][9] ), .B(n10729), .Y(n1228) );
  INVX1 U8076 ( .A(n1228), .Y(n6099) );
  AND2X1 U8077 ( .A(\RF[15][63] ), .B(n10731), .Y(n1216) );
  INVX1 U8078 ( .A(n1216), .Y(n6100) );
  AND2X1 U8079 ( .A(\RF[15][34] ), .B(n10731), .Y(n1187) );
  INVX1 U8080 ( .A(n1187), .Y(n6101) );
  AND2X1 U8081 ( .A(\RF[15][22] ), .B(n10732), .Y(n1175) );
  INVX1 U8082 ( .A(n1175), .Y(n6102) );
  AND2X1 U8083 ( .A(\RF[15][10] ), .B(n10731), .Y(n1163) );
  INVX1 U8084 ( .A(n1163), .Y(n6103) );
  AND2X1 U8085 ( .A(\RF[16][43] ), .B(n10733), .Y(n1131) );
  INVX1 U8086 ( .A(n1131), .Y(n6104) );
  AND2X1 U8087 ( .A(\RF[16][31] ), .B(n10733), .Y(n1119) );
  INVX1 U8088 ( .A(n1119), .Y(n6105) );
  AND2X1 U8089 ( .A(\RF[16][19] ), .B(n10734), .Y(n1107) );
  INVX1 U8090 ( .A(n1107), .Y(n6106) );
  AND2X1 U8091 ( .A(\RF[16][7] ), .B(n10733), .Y(n1095) );
  INVX1 U8092 ( .A(n1095), .Y(n6107) );
  AND2X1 U8093 ( .A(\RF[17][47] ), .B(n10735), .Y(n1070) );
  INVX1 U8094 ( .A(n1070), .Y(n6108) );
  AND2X1 U8095 ( .A(\RF[17][25] ), .B(n10735), .Y(n1048) );
  INVX1 U8096 ( .A(n1048), .Y(n6109) );
  AND2X1 U8097 ( .A(\RF[17][20] ), .B(n10736), .Y(n1043) );
  INVX1 U8098 ( .A(n1043), .Y(n6110) );
  AND2X1 U8099 ( .A(\RF[17][8] ), .B(n10735), .Y(n1031) );
  INVX1 U8100 ( .A(n1031), .Y(n6111) );
  AND2X1 U8101 ( .A(\RF[18][41] ), .B(n10737), .Y(n999) );
  INVX1 U8102 ( .A(n999), .Y(n6112) );
  AND2X1 U8103 ( .A(\RF[18][29] ), .B(n10738), .Y(n987) );
  INVX1 U8104 ( .A(n987), .Y(n6113) );
  AND2X1 U8105 ( .A(\RF[18][17] ), .B(n10737), .Y(n975) );
  INVX1 U8106 ( .A(n975), .Y(n6114) );
  AND2X1 U8107 ( .A(\RF[18][5] ), .B(n10737), .Y(n963) );
  INVX1 U8108 ( .A(n963), .Y(n6115) );
  AND2X1 U8109 ( .A(\RF[19][38] ), .B(n10740), .Y(n931) );
  INVX1 U8110 ( .A(n931), .Y(n6116) );
  AND2X1 U8111 ( .A(\RF[19][30] ), .B(n10739), .Y(n923) );
  INVX1 U8112 ( .A(n923), .Y(n6117) );
  AND2X1 U8113 ( .A(\RF[19][18] ), .B(n10739), .Y(n911) );
  INVX1 U8114 ( .A(n911), .Y(n6118) );
  AND2X1 U8115 ( .A(\RF[19][6] ), .B(n10739), .Y(n899) );
  INVX1 U8116 ( .A(n899), .Y(n6119) );
  AND2X1 U8117 ( .A(\RF[20][39] ), .B(n10741), .Y(n867) );
  INVX1 U8118 ( .A(n867), .Y(n6120) );
  AND2X1 U8119 ( .A(\RF[20][27] ), .B(n10742), .Y(n855) );
  INVX1 U8120 ( .A(n855), .Y(n6121) );
  AND2X1 U8121 ( .A(\RF[20][15] ), .B(n10741), .Y(n843) );
  INVX1 U8122 ( .A(n843), .Y(n6122) );
  AND2X1 U8123 ( .A(\RF[20][3] ), .B(n10741), .Y(n831) );
  INVX1 U8124 ( .A(n831), .Y(n6123) );
  AND2X1 U8125 ( .A(\RF[21][40] ), .B(n10743), .Y(n803) );
  INVX1 U8126 ( .A(n803), .Y(n6124) );
  AND2X1 U8127 ( .A(\RF[21][28] ), .B(n10744), .Y(n791) );
  INVX1 U8128 ( .A(n791), .Y(n6125) );
  AND2X1 U8129 ( .A(\RF[21][16] ), .B(n10743), .Y(n779) );
  INVX1 U8130 ( .A(n779), .Y(n6126) );
  AND2X1 U8131 ( .A(\RF[21][4] ), .B(n10743), .Y(n767) );
  INVX1 U8132 ( .A(n767), .Y(n6127) );
  AND2X1 U8133 ( .A(\RF[22][45] ), .B(n10746), .Y(n743) );
  INVX1 U8134 ( .A(n743), .Y(n6128) );
  AND2X1 U8135 ( .A(\RF[22][32] ), .B(n10745), .Y(n730) );
  INVX1 U8136 ( .A(n730), .Y(n6129) );
  AND2X1 U8137 ( .A(\RF[22][13] ), .B(n10745), .Y(n711) );
  INVX1 U8138 ( .A(n711), .Y(n6130) );
  AND2X1 U8139 ( .A(\RF[22][1] ), .B(n10745), .Y(n699) );
  INVX1 U8140 ( .A(n699), .Y(n6131) );
  AND2X1 U8141 ( .A(\RF[22][0] ), .B(n10745), .Y(n698) );
  INVX1 U8142 ( .A(n698), .Y(n6132) );
  AND2X1 U8143 ( .A(\RF[23][37] ), .B(n10747), .Y(n669) );
  INVX1 U8144 ( .A(n669), .Y(n6133) );
  AND2X1 U8145 ( .A(\RF[23][26] ), .B(n10748), .Y(n658) );
  INVX1 U8146 ( .A(n658), .Y(n6134) );
  AND2X1 U8147 ( .A(\RF[23][14] ), .B(n10747), .Y(n646) );
  INVX1 U8148 ( .A(n646), .Y(n6135) );
  AND2X1 U8149 ( .A(\RF[23][2] ), .B(n10747), .Y(n634) );
  INVX1 U8150 ( .A(n634), .Y(n6136) );
  AND2X1 U8151 ( .A(\RF[24][43] ), .B(n10749), .Y(n608) );
  INVX1 U8152 ( .A(n608), .Y(n6137) );
  AND2X1 U8153 ( .A(\RF[24][31] ), .B(n10749), .Y(n596) );
  INVX1 U8154 ( .A(n596), .Y(n6138) );
  AND2X1 U8155 ( .A(\RF[24][19] ), .B(n10750), .Y(n584) );
  INVX1 U8156 ( .A(n584), .Y(n6139) );
  AND2X1 U8157 ( .A(\RF[24][7] ), .B(n10749), .Y(n572) );
  INVX1 U8158 ( .A(n572), .Y(n6140) );
  AND2X1 U8159 ( .A(\RF[25][47] ), .B(n10751), .Y(n546) );
  INVX1 U8160 ( .A(n546), .Y(n6141) );
  AND2X1 U8161 ( .A(\RF[25][25] ), .B(n10751), .Y(n524) );
  INVX1 U8162 ( .A(n524), .Y(n6142) );
  AND2X1 U8163 ( .A(\RF[25][20] ), .B(n10752), .Y(n519) );
  INVX1 U8164 ( .A(n519), .Y(n6143) );
  AND2X1 U8165 ( .A(\RF[25][8] ), .B(n10751), .Y(n507) );
  INVX1 U8166 ( .A(n507), .Y(n6144) );
  AND2X1 U8167 ( .A(\RF[26][41] ), .B(n10753), .Y(n474) );
  INVX1 U8168 ( .A(n474), .Y(n6145) );
  AND2X1 U8169 ( .A(\RF[26][29] ), .B(n10754), .Y(n462) );
  INVX1 U8170 ( .A(n462), .Y(n6146) );
  AND2X1 U8171 ( .A(\RF[26][17] ), .B(n10753), .Y(n450) );
  INVX1 U8172 ( .A(n450), .Y(n6147) );
  AND2X1 U8173 ( .A(\RF[26][5] ), .B(n10753), .Y(n438) );
  INVX1 U8174 ( .A(n438), .Y(n6148) );
  AND2X1 U8175 ( .A(\RF[27][38] ), .B(n10756), .Y(n405) );
  INVX1 U8176 ( .A(n405), .Y(n6149) );
  AND2X1 U8177 ( .A(\RF[27][30] ), .B(n10755), .Y(n397) );
  INVX1 U8178 ( .A(n397), .Y(n6150) );
  AND2X1 U8179 ( .A(\RF[27][18] ), .B(n10755), .Y(n385) );
  INVX1 U8180 ( .A(n385), .Y(n6151) );
  AND2X1 U8181 ( .A(\RF[27][6] ), .B(n10755), .Y(n373) );
  INVX1 U8182 ( .A(n373), .Y(n6152) );
  AND2X1 U8183 ( .A(\RF[28][39] ), .B(n10757), .Y(n340) );
  INVX1 U8184 ( .A(n340), .Y(n6153) );
  AND2X1 U8185 ( .A(\RF[28][27] ), .B(n10758), .Y(n328) );
  INVX1 U8186 ( .A(n328), .Y(n6154) );
  AND2X1 U8187 ( .A(\RF[28][15] ), .B(n10757), .Y(n316) );
  INVX1 U8188 ( .A(n316), .Y(n6155) );
  AND2X1 U8189 ( .A(\RF[28][3] ), .B(n10757), .Y(n304) );
  INVX1 U8190 ( .A(n304), .Y(n6156) );
  AND2X1 U8191 ( .A(\RF[29][40] ), .B(n10759), .Y(n275) );
  INVX1 U8192 ( .A(n275), .Y(n6157) );
  AND2X1 U8193 ( .A(\RF[29][28] ), .B(n10760), .Y(n263) );
  INVX1 U8194 ( .A(n263), .Y(n6158) );
  AND2X1 U8195 ( .A(\RF[29][16] ), .B(n10759), .Y(n251) );
  INVX1 U8196 ( .A(n251), .Y(n6159) );
  AND2X1 U8197 ( .A(\RF[29][4] ), .B(n10759), .Y(n239) );
  INVX1 U8198 ( .A(n239), .Y(n6160) );
  AND2X1 U8199 ( .A(\RF[30][45] ), .B(n10762), .Y(n214) );
  INVX1 U8200 ( .A(n214), .Y(n6161) );
  AND2X1 U8201 ( .A(\RF[30][32] ), .B(n10761), .Y(n201) );
  INVX1 U8202 ( .A(n201), .Y(n6162) );
  AND2X1 U8203 ( .A(\RF[30][13] ), .B(n10761), .Y(n182) );
  INVX1 U8204 ( .A(n182), .Y(n6163) );
  AND2X1 U8205 ( .A(\RF[30][1] ), .B(n10761), .Y(n170) );
  INVX1 U8206 ( .A(n170), .Y(n6164) );
  AND2X1 U8207 ( .A(\RF[30][0] ), .B(n10761), .Y(n169) );
  INVX1 U8208 ( .A(n169), .Y(n6165) );
  AND2X1 U8209 ( .A(\RF[31][37] ), .B(n10763), .Y(n113) );
  INVX1 U8210 ( .A(n113), .Y(n6166) );
  AND2X1 U8211 ( .A(\RF[31][26] ), .B(n10764), .Y(n91) );
  INVX1 U8212 ( .A(n91), .Y(n6167) );
  AND2X1 U8213 ( .A(\RF[31][14] ), .B(n10763), .Y(n67) );
  INVX1 U8214 ( .A(n67), .Y(n6168) );
  AND2X1 U8215 ( .A(\RF[31][2] ), .B(n10763), .Y(n43) );
  INVX1 U8216 ( .A(n43), .Y(n6169) );
  BUFX2 U8217 ( .A(n1218), .Y(n6170) );
  AND2X1 U8218 ( .A(\RF[0][59] ), .B(n10702), .Y(n2189) );
  INVX1 U8219 ( .A(n2189), .Y(n6171) );
  AND2X1 U8220 ( .A(\RF[0][42] ), .B(n10702), .Y(n2172) );
  INVX1 U8221 ( .A(n2172), .Y(n6172) );
  AND2X1 U8222 ( .A(\RF[0][36] ), .B(n10702), .Y(n2166) );
  INVX1 U8223 ( .A(n2166), .Y(n6173) );
  AND2X1 U8224 ( .A(\RF[0][12] ), .B(n10702), .Y(n2142) );
  INVX1 U8225 ( .A(n2142), .Y(n6174) );
  AND2X1 U8226 ( .A(\RF[1][56] ), .B(n10704), .Y(n2121) );
  INVX1 U8227 ( .A(n2121), .Y(n6175) );
  AND2X1 U8228 ( .A(\RF[1][35] ), .B(n10704), .Y(n2100) );
  INVX1 U8229 ( .A(n2100), .Y(n6176) );
  AND2X1 U8230 ( .A(\RF[1][23] ), .B(n10704), .Y(n2088) );
  INVX1 U8231 ( .A(n2088), .Y(n6177) );
  AND2X1 U8232 ( .A(\RF[1][11] ), .B(n10704), .Y(n2076) );
  INVX1 U8233 ( .A(n2076), .Y(n6178) );
  AND2X1 U8234 ( .A(\RF[2][63] ), .B(n10705), .Y(n2063) );
  INVX1 U8235 ( .A(n2063), .Y(n6179) );
  AND2X1 U8236 ( .A(\RF[2][34] ), .B(n10706), .Y(n2034) );
  INVX1 U8237 ( .A(n2034), .Y(n6180) );
  AND2X1 U8238 ( .A(\RF[2][22] ), .B(n10706), .Y(n2022) );
  INVX1 U8239 ( .A(n2022), .Y(n6181) );
  AND2X1 U8240 ( .A(\RF[2][10] ), .B(n10705), .Y(n2010) );
  INVX1 U8241 ( .A(n2010), .Y(n6182) );
  AND2X1 U8242 ( .A(\RF[3][44] ), .B(n10708), .Y(n1979) );
  INVX1 U8243 ( .A(n1979), .Y(n6183) );
  AND2X1 U8244 ( .A(\RF[3][33] ), .B(n10708), .Y(n1968) );
  INVX1 U8245 ( .A(n1968), .Y(n6184) );
  AND2X1 U8246 ( .A(\RF[3][21] ), .B(n10708), .Y(n1956) );
  INVX1 U8247 ( .A(n1956), .Y(n6185) );
  AND2X1 U8248 ( .A(\RF[3][9] ), .B(n10708), .Y(n1944) );
  INVX1 U8249 ( .A(n1944), .Y(n6186) );
  AND2X1 U8250 ( .A(\RF[4][47] ), .B(n10710), .Y(n1917) );
  INVX1 U8251 ( .A(n1917), .Y(n6187) );
  AND2X1 U8252 ( .A(\RF[4][25] ), .B(n10710), .Y(n1895) );
  INVX1 U8253 ( .A(n1895), .Y(n6188) );
  AND2X1 U8254 ( .A(\RF[4][20] ), .B(n10710), .Y(n1890) );
  INVX1 U8255 ( .A(n1890), .Y(n6189) );
  AND2X1 U8256 ( .A(\RF[4][8] ), .B(n10710), .Y(n1878) );
  INVX1 U8257 ( .A(n1878), .Y(n6190) );
  AND2X1 U8258 ( .A(\RF[5][43] ), .B(n10712), .Y(n1848) );
  INVX1 U8259 ( .A(n1848), .Y(n6191) );
  AND2X1 U8260 ( .A(\RF[5][31] ), .B(n10712), .Y(n1836) );
  INVX1 U8261 ( .A(n1836), .Y(n6192) );
  AND2X1 U8262 ( .A(\RF[5][19] ), .B(n10712), .Y(n1824) );
  INVX1 U8263 ( .A(n1824), .Y(n6193) );
  AND2X1 U8264 ( .A(\RF[5][7] ), .B(n10711), .Y(n1812) );
  INVX1 U8265 ( .A(n1812), .Y(n6194) );
  AND2X1 U8266 ( .A(\RF[6][38] ), .B(n10714), .Y(n1778) );
  INVX1 U8267 ( .A(n1778), .Y(n6195) );
  AND2X1 U8268 ( .A(\RF[6][30] ), .B(n10714), .Y(n1770) );
  INVX1 U8269 ( .A(n1770), .Y(n6196) );
  AND2X1 U8270 ( .A(\RF[6][18] ), .B(n10714), .Y(n1758) );
  INVX1 U8271 ( .A(n1758), .Y(n6197) );
  AND2X1 U8272 ( .A(\RF[6][6] ), .B(n10713), .Y(n1746) );
  INVX1 U8273 ( .A(n1746), .Y(n6198) );
  AND2X1 U8274 ( .A(\RF[7][41] ), .B(n10716), .Y(n1715) );
  INVX1 U8275 ( .A(n1715), .Y(n6199) );
  AND2X1 U8276 ( .A(\RF[7][29] ), .B(n10716), .Y(n1703) );
  INVX1 U8277 ( .A(n1703), .Y(n6200) );
  AND2X1 U8278 ( .A(\RF[7][17] ), .B(n10716), .Y(n1691) );
  INVX1 U8279 ( .A(n1691), .Y(n6201) );
  AND2X1 U8280 ( .A(\RF[7][5] ), .B(n10715), .Y(n1679) );
  INVX1 U8281 ( .A(n1679), .Y(n6202) );
  AND2X1 U8282 ( .A(\RF[8][40] ), .B(n10718), .Y(n1649) );
  INVX1 U8283 ( .A(n1649), .Y(n6203) );
  AND2X1 U8284 ( .A(\RF[8][28] ), .B(n10718), .Y(n1637) );
  INVX1 U8285 ( .A(n1637), .Y(n6204) );
  AND2X1 U8286 ( .A(\RF[8][16] ), .B(n10718), .Y(n1625) );
  INVX1 U8287 ( .A(n1625), .Y(n6205) );
  AND2X1 U8288 ( .A(\RF[8][4] ), .B(n10717), .Y(n1613) );
  INVX1 U8289 ( .A(n1613), .Y(n6206) );
  AND2X1 U8290 ( .A(\RF[9][39] ), .B(n10720), .Y(n1583) );
  INVX1 U8291 ( .A(n1583), .Y(n6207) );
  AND2X1 U8292 ( .A(\RF[9][27] ), .B(n10720), .Y(n1571) );
  INVX1 U8293 ( .A(n1571), .Y(n6208) );
  AND2X1 U8294 ( .A(\RF[9][15] ), .B(n10720), .Y(n1559) );
  INVX1 U8295 ( .A(n1559), .Y(n6209) );
  AND2X1 U8296 ( .A(\RF[9][3] ), .B(n10719), .Y(n1547) );
  INVX1 U8297 ( .A(n1547), .Y(n6210) );
  AND2X1 U8298 ( .A(\RF[10][37] ), .B(n10722), .Y(n1516) );
  INVX1 U8299 ( .A(n1516), .Y(n6211) );
  AND2X1 U8300 ( .A(\RF[10][26] ), .B(n10722), .Y(n1505) );
  INVX1 U8301 ( .A(n1505), .Y(n6212) );
  AND2X1 U8302 ( .A(\RF[10][14] ), .B(n10722), .Y(n1493) );
  INVX1 U8303 ( .A(n1493), .Y(n6213) );
  AND2X1 U8304 ( .A(\RF[10][2] ), .B(n10721), .Y(n1481) );
  INVX1 U8305 ( .A(n1481), .Y(n6214) );
  AND2X1 U8306 ( .A(\RF[11][45] ), .B(n10724), .Y(n1459) );
  INVX1 U8307 ( .A(n1459), .Y(n6215) );
  AND2X1 U8308 ( .A(\RF[11][32] ), .B(n10724), .Y(n1446) );
  INVX1 U8309 ( .A(n1446), .Y(n6216) );
  AND2X1 U8310 ( .A(\RF[11][13] ), .B(n10724), .Y(n1427) );
  INVX1 U8311 ( .A(n1427), .Y(n6217) );
  AND2X1 U8312 ( .A(\RF[11][1] ), .B(n10723), .Y(n1415) );
  INVX1 U8313 ( .A(n1415), .Y(n6218) );
  AND2X1 U8314 ( .A(\RF[11][0] ), .B(n10723), .Y(n1414) );
  INVX1 U8315 ( .A(n1414), .Y(n6219) );
  AND2X1 U8316 ( .A(\RF[12][59] ), .B(n10726), .Y(n1408) );
  INVX1 U8317 ( .A(n1408), .Y(n6220) );
  AND2X1 U8318 ( .A(\RF[12][42] ), .B(n10726), .Y(n1391) );
  INVX1 U8319 ( .A(n1391), .Y(n6221) );
  AND2X1 U8320 ( .A(\RF[12][36] ), .B(n10726), .Y(n1385) );
  INVX1 U8321 ( .A(n1385), .Y(n6222) );
  AND2X1 U8322 ( .A(\RF[12][12] ), .B(n10726), .Y(n1361) );
  INVX1 U8323 ( .A(n1361), .Y(n6223) );
  AND2X1 U8324 ( .A(\RF[13][56] ), .B(n10728), .Y(n1340) );
  INVX1 U8325 ( .A(n1340), .Y(n6224) );
  AND2X1 U8326 ( .A(\RF[13][35] ), .B(n10728), .Y(n1319) );
  INVX1 U8327 ( .A(n1319), .Y(n6225) );
  AND2X1 U8328 ( .A(\RF[13][23] ), .B(n10728), .Y(n1307) );
  INVX1 U8329 ( .A(n1307), .Y(n6226) );
  AND2X1 U8330 ( .A(\RF[13][11] ), .B(n10728), .Y(n1295) );
  INVX1 U8331 ( .A(n1295), .Y(n6227) );
  AND2X1 U8332 ( .A(\RF[14][63] ), .B(n10729), .Y(n1282) );
  INVX1 U8333 ( .A(n1282), .Y(n6228) );
  AND2X1 U8334 ( .A(\RF[14][34] ), .B(n10730), .Y(n1253) );
  INVX1 U8335 ( .A(n1253), .Y(n6229) );
  AND2X1 U8336 ( .A(\RF[14][22] ), .B(n10730), .Y(n1241) );
  INVX1 U8337 ( .A(n1241), .Y(n6230) );
  AND2X1 U8338 ( .A(\RF[14][10] ), .B(n10729), .Y(n1229) );
  INVX1 U8339 ( .A(n1229), .Y(n6231) );
  AND2X1 U8340 ( .A(\RF[15][44] ), .B(n10732), .Y(n1197) );
  INVX1 U8341 ( .A(n1197), .Y(n6232) );
  AND2X1 U8342 ( .A(\RF[15][33] ), .B(n10732), .Y(n1186) );
  INVX1 U8343 ( .A(n1186), .Y(n6233) );
  AND2X1 U8344 ( .A(\RF[15][21] ), .B(n10732), .Y(n1174) );
  INVX1 U8345 ( .A(n1174), .Y(n6234) );
  AND2X1 U8346 ( .A(\RF[15][9] ), .B(n10732), .Y(n1162) );
  INVX1 U8347 ( .A(n1162), .Y(n6235) );
  AND2X1 U8348 ( .A(\RF[16][47] ), .B(n10734), .Y(n1135) );
  INVX1 U8349 ( .A(n1135), .Y(n6236) );
  AND2X1 U8350 ( .A(\RF[16][25] ), .B(n10734), .Y(n1113) );
  INVX1 U8351 ( .A(n1113), .Y(n6237) );
  AND2X1 U8352 ( .A(\RF[16][20] ), .B(n10734), .Y(n1108) );
  INVX1 U8353 ( .A(n1108), .Y(n6238) );
  AND2X1 U8354 ( .A(\RF[16][8] ), .B(n10734), .Y(n1096) );
  INVX1 U8355 ( .A(n1096), .Y(n6239) );
  AND2X1 U8356 ( .A(\RF[17][43] ), .B(n10736), .Y(n1066) );
  INVX1 U8357 ( .A(n1066), .Y(n6240) );
  AND2X1 U8358 ( .A(\RF[17][31] ), .B(n10736), .Y(n1054) );
  INVX1 U8359 ( .A(n1054), .Y(n6241) );
  AND2X1 U8360 ( .A(\RF[17][19] ), .B(n10736), .Y(n1042) );
  INVX1 U8361 ( .A(n1042), .Y(n6242) );
  AND2X1 U8362 ( .A(\RF[17][7] ), .B(n10735), .Y(n1030) );
  INVX1 U8363 ( .A(n1030), .Y(n6243) );
  AND2X1 U8364 ( .A(\RF[18][38] ), .B(n10738), .Y(n996) );
  INVX1 U8365 ( .A(n996), .Y(n6244) );
  AND2X1 U8366 ( .A(\RF[18][30] ), .B(n10738), .Y(n988) );
  INVX1 U8367 ( .A(n988), .Y(n6245) );
  AND2X1 U8368 ( .A(\RF[18][18] ), .B(n10738), .Y(n976) );
  INVX1 U8369 ( .A(n976), .Y(n6246) );
  AND2X1 U8370 ( .A(\RF[18][6] ), .B(n10737), .Y(n964) );
  INVX1 U8371 ( .A(n964), .Y(n6247) );
  AND2X1 U8372 ( .A(\RF[19][41] ), .B(n10740), .Y(n934) );
  INVX1 U8373 ( .A(n934), .Y(n6248) );
  AND2X1 U8374 ( .A(\RF[19][29] ), .B(n10740), .Y(n922) );
  INVX1 U8375 ( .A(n922), .Y(n6249) );
  AND2X1 U8376 ( .A(\RF[19][17] ), .B(n10740), .Y(n910) );
  INVX1 U8377 ( .A(n910), .Y(n6250) );
  AND2X1 U8378 ( .A(\RF[19][5] ), .B(n10739), .Y(n898) );
  INVX1 U8379 ( .A(n898), .Y(n6251) );
  AND2X1 U8380 ( .A(\RF[20][40] ), .B(n10742), .Y(n868) );
  INVX1 U8381 ( .A(n868), .Y(n6252) );
  AND2X1 U8382 ( .A(\RF[20][28] ), .B(n10742), .Y(n856) );
  INVX1 U8383 ( .A(n856), .Y(n6253) );
  AND2X1 U8384 ( .A(\RF[20][16] ), .B(n10742), .Y(n844) );
  INVX1 U8385 ( .A(n844), .Y(n6254) );
  AND2X1 U8386 ( .A(\RF[20][4] ), .B(n10741), .Y(n832) );
  INVX1 U8387 ( .A(n832), .Y(n6255) );
  AND2X1 U8388 ( .A(\RF[21][39] ), .B(n10744), .Y(n802) );
  INVX1 U8389 ( .A(n802), .Y(n6256) );
  AND2X1 U8390 ( .A(\RF[21][27] ), .B(n10744), .Y(n790) );
  INVX1 U8391 ( .A(n790), .Y(n6257) );
  AND2X1 U8392 ( .A(\RF[21][15] ), .B(n10744), .Y(n778) );
  INVX1 U8393 ( .A(n778), .Y(n6258) );
  AND2X1 U8394 ( .A(\RF[21][3] ), .B(n10743), .Y(n766) );
  INVX1 U8395 ( .A(n766), .Y(n6259) );
  AND2X1 U8396 ( .A(\RF[22][37] ), .B(n10746), .Y(n735) );
  INVX1 U8397 ( .A(n735), .Y(n6260) );
  AND2X1 U8398 ( .A(\RF[22][26] ), .B(n10746), .Y(n724) );
  INVX1 U8399 ( .A(n724), .Y(n6261) );
  AND2X1 U8400 ( .A(\RF[22][14] ), .B(n10746), .Y(n712) );
  INVX1 U8401 ( .A(n712), .Y(n6262) );
  AND2X1 U8402 ( .A(\RF[22][2] ), .B(n10745), .Y(n700) );
  INVX1 U8403 ( .A(n700), .Y(n6263) );
  AND2X1 U8404 ( .A(\RF[23][45] ), .B(n10748), .Y(n677) );
  INVX1 U8405 ( .A(n677), .Y(n6264) );
  AND2X1 U8406 ( .A(\RF[23][32] ), .B(n10748), .Y(n664) );
  INVX1 U8407 ( .A(n664), .Y(n6265) );
  AND2X1 U8408 ( .A(\RF[23][13] ), .B(n10748), .Y(n645) );
  INVX1 U8409 ( .A(n645), .Y(n6266) );
  AND2X1 U8410 ( .A(\RF[23][1] ), .B(n10747), .Y(n633) );
  INVX1 U8411 ( .A(n633), .Y(n6267) );
  AND2X1 U8412 ( .A(\RF[23][0] ), .B(n10747), .Y(n632) );
  INVX1 U8413 ( .A(n632), .Y(n6268) );
  AND2X1 U8414 ( .A(\RF[24][47] ), .B(n10750), .Y(n612) );
  INVX1 U8415 ( .A(n612), .Y(n6269) );
  AND2X1 U8416 ( .A(\RF[24][25] ), .B(n10750), .Y(n590) );
  INVX1 U8417 ( .A(n590), .Y(n6270) );
  AND2X1 U8418 ( .A(\RF[24][20] ), .B(n10750), .Y(n585) );
  INVX1 U8419 ( .A(n585), .Y(n6271) );
  AND2X1 U8420 ( .A(\RF[24][8] ), .B(n10750), .Y(n573) );
  INVX1 U8421 ( .A(n573), .Y(n6272) );
  AND2X1 U8422 ( .A(\RF[25][43] ), .B(n10752), .Y(n542) );
  INVX1 U8423 ( .A(n542), .Y(n6273) );
  AND2X1 U8424 ( .A(\RF[25][31] ), .B(n10752), .Y(n530) );
  INVX1 U8425 ( .A(n530), .Y(n6274) );
  AND2X1 U8426 ( .A(\RF[25][19] ), .B(n10752), .Y(n518) );
  INVX1 U8427 ( .A(n518), .Y(n6275) );
  AND2X1 U8428 ( .A(\RF[25][7] ), .B(n10751), .Y(n506) );
  INVX1 U8429 ( .A(n506), .Y(n6276) );
  AND2X1 U8430 ( .A(\RF[26][38] ), .B(n10754), .Y(n471) );
  INVX1 U8431 ( .A(n471), .Y(n6277) );
  AND2X1 U8432 ( .A(\RF[26][30] ), .B(n10754), .Y(n463) );
  INVX1 U8433 ( .A(n463), .Y(n6278) );
  AND2X1 U8434 ( .A(\RF[26][18] ), .B(n10754), .Y(n451) );
  INVX1 U8435 ( .A(n451), .Y(n6279) );
  AND2X1 U8436 ( .A(\RF[26][6] ), .B(n10753), .Y(n439) );
  INVX1 U8437 ( .A(n439), .Y(n6280) );
  AND2X1 U8438 ( .A(\RF[27][41] ), .B(n10756), .Y(n408) );
  INVX1 U8439 ( .A(n408), .Y(n6281) );
  AND2X1 U8440 ( .A(\RF[27][29] ), .B(n10756), .Y(n396) );
  INVX1 U8441 ( .A(n396), .Y(n6282) );
  AND2X1 U8442 ( .A(\RF[27][17] ), .B(n10756), .Y(n384) );
  INVX1 U8443 ( .A(n384), .Y(n6283) );
  AND2X1 U8444 ( .A(\RF[27][5] ), .B(n10755), .Y(n372) );
  INVX1 U8445 ( .A(n372), .Y(n6284) );
  AND2X1 U8446 ( .A(\RF[28][40] ), .B(n10758), .Y(n341) );
  INVX1 U8447 ( .A(n341), .Y(n6285) );
  AND2X1 U8448 ( .A(\RF[28][28] ), .B(n10758), .Y(n329) );
  INVX1 U8449 ( .A(n329), .Y(n6286) );
  AND2X1 U8450 ( .A(\RF[28][16] ), .B(n10758), .Y(n317) );
  INVX1 U8451 ( .A(n317), .Y(n6287) );
  AND2X1 U8452 ( .A(\RF[28][4] ), .B(n10757), .Y(n305) );
  INVX1 U8453 ( .A(n305), .Y(n6288) );
  AND2X1 U8454 ( .A(\RF[29][39] ), .B(n10760), .Y(n274) );
  INVX1 U8455 ( .A(n274), .Y(n6289) );
  AND2X1 U8456 ( .A(\RF[29][27] ), .B(n10760), .Y(n262) );
  INVX1 U8457 ( .A(n262), .Y(n6290) );
  AND2X1 U8458 ( .A(\RF[29][15] ), .B(n10760), .Y(n250) );
  INVX1 U8459 ( .A(n250), .Y(n6291) );
  AND2X1 U8460 ( .A(\RF[29][3] ), .B(n10759), .Y(n238) );
  INVX1 U8461 ( .A(n238), .Y(n6292) );
  AND2X1 U8462 ( .A(\RF[30][37] ), .B(n10762), .Y(n206) );
  INVX1 U8463 ( .A(n206), .Y(n6293) );
  AND2X1 U8464 ( .A(\RF[30][26] ), .B(n10762), .Y(n195) );
  INVX1 U8465 ( .A(n195), .Y(n6294) );
  AND2X1 U8466 ( .A(\RF[30][14] ), .B(n10762), .Y(n183) );
  INVX1 U8467 ( .A(n183), .Y(n6295) );
  AND2X1 U8468 ( .A(\RF[30][2] ), .B(n10761), .Y(n171) );
  INVX1 U8469 ( .A(n171), .Y(n6296) );
  AND2X1 U8470 ( .A(\RF[31][45] ), .B(n10764), .Y(n129) );
  INVX1 U8471 ( .A(n129), .Y(n6297) );
  AND2X1 U8472 ( .A(\RF[31][32] ), .B(n10764), .Y(n103) );
  INVX1 U8473 ( .A(n103), .Y(n6298) );
  AND2X1 U8474 ( .A(\RF[31][13] ), .B(n10764), .Y(n65) );
  INVX1 U8475 ( .A(n65), .Y(n6299) );
  AND2X1 U8476 ( .A(\RF[31][1] ), .B(n10763), .Y(n41) );
  INVX1 U8477 ( .A(n41), .Y(n6300) );
  AND2X1 U8478 ( .A(\RF[31][0] ), .B(n10763), .Y(n39) );
  INVX1 U8479 ( .A(n39), .Y(n6301) );
  BUFX2 U8480 ( .A(n697), .Y(n6302) );
  INVX1 U8481 ( .A(n10534), .Y(n10547) );
  INVX1 U8482 ( .A(n10534), .Y(n10548) );
  INVX1 U8483 ( .A(n10534), .Y(n10549) );
  INVX1 U8484 ( .A(n10533), .Y(n10550) );
  INVX1 U8485 ( .A(n10533), .Y(n10551) );
  INVX1 U8486 ( .A(n10533), .Y(n10552) );
  INVX1 U8487 ( .A(n10532), .Y(n10553) );
  INVX1 U8488 ( .A(n10532), .Y(n10554) );
  INVX1 U8489 ( .A(n10532), .Y(n10555) );
  INVX1 U8490 ( .A(n10531), .Y(n10556) );
  INVX1 U8491 ( .A(n10531), .Y(n10557) );
  INVX1 U8492 ( .A(n10531), .Y(n10558) );
  INVX1 U8493 ( .A(n10530), .Y(n10559) );
  INVX1 U8494 ( .A(n10530), .Y(n10560) );
  INVX1 U8495 ( .A(n10530), .Y(n10561) );
  INVX1 U8496 ( .A(n10529), .Y(n10562) );
  INVX1 U8497 ( .A(n10529), .Y(n10563) );
  INVX1 U8498 ( .A(n10529), .Y(n10564) );
  INVX1 U8499 ( .A(n10528), .Y(n10565) );
  INVX1 U8500 ( .A(n10528), .Y(n10566) );
  INVX1 U8501 ( .A(n10528), .Y(n10567) );
  INVX1 U8502 ( .A(n10527), .Y(n10568) );
  INVX1 U8503 ( .A(n10527), .Y(n10569) );
  INVX1 U8504 ( .A(n10527), .Y(n10570) );
  INVX1 U8505 ( .A(n10626), .Y(n10571) );
  INVX1 U8506 ( .A(n10537), .Y(n10572) );
  INVX1 U8507 ( .A(n10536), .Y(n10573) );
  INVX1 U8508 ( .A(n10526), .Y(n10574) );
  INVX1 U8509 ( .A(n10526), .Y(n10575) );
  INVX1 U8510 ( .A(n10526), .Y(n10576) );
  INVX1 U8511 ( .A(n10525), .Y(n10577) );
  INVX1 U8512 ( .A(n10525), .Y(n10578) );
  INVX1 U8513 ( .A(n10525), .Y(n10579) );
  INVX1 U8514 ( .A(n10524), .Y(n10580) );
  INVX1 U8515 ( .A(n10524), .Y(n10581) );
  INVX1 U8516 ( .A(n10524), .Y(n10582) );
  INVX1 U8517 ( .A(n10523), .Y(n10583) );
  INVX1 U8518 ( .A(n10523), .Y(n10584) );
  INVX1 U8519 ( .A(n10523), .Y(n10585) );
  INVX1 U8520 ( .A(n10522), .Y(n10586) );
  INVX1 U8521 ( .A(n10522), .Y(n10587) );
  INVX1 U8522 ( .A(n10522), .Y(n10588) );
  INVX1 U8523 ( .A(n10521), .Y(n10589) );
  INVX1 U8524 ( .A(n10521), .Y(n10590) );
  INVX1 U8525 ( .A(n10521), .Y(n10591) );
  INVX1 U8526 ( .A(n10523), .Y(n10592) );
  INVX1 U8527 ( .A(n10522), .Y(n10593) );
  INVX1 U8528 ( .A(n10521), .Y(n10594) );
  INVX1 U8529 ( .A(n10628), .Y(n10595) );
  INVX1 U8530 ( .A(n10525), .Y(n10596) );
  INVX1 U8531 ( .A(n10524), .Y(n10597) );
  INVX1 U8532 ( .A(n10531), .Y(n10598) );
  INVX1 U8533 ( .A(n10530), .Y(n10599) );
  INVX1 U8534 ( .A(n10529), .Y(n10600) );
  INVX1 U8535 ( .A(n8367), .Y(n8380) );
  INVX1 U8536 ( .A(n8367), .Y(n8381) );
  INVX1 U8537 ( .A(n8367), .Y(n8382) );
  INVX1 U8538 ( .A(n8366), .Y(n8383) );
  INVX1 U8539 ( .A(n8366), .Y(n8384) );
  INVX1 U8540 ( .A(n8366), .Y(n8385) );
  INVX1 U8541 ( .A(n8365), .Y(n8386) );
  INVX1 U8542 ( .A(n8365), .Y(n8387) );
  INVX1 U8543 ( .A(n8365), .Y(n8388) );
  INVX1 U8544 ( .A(n8364), .Y(n8389) );
  INVX1 U8545 ( .A(n8364), .Y(n8390) );
  INVX1 U8546 ( .A(n8364), .Y(n8391) );
  INVX1 U8547 ( .A(n8363), .Y(n8392) );
  INVX1 U8548 ( .A(n8363), .Y(n8393) );
  INVX1 U8549 ( .A(n8363), .Y(n8394) );
  INVX1 U8550 ( .A(n8362), .Y(n8395) );
  INVX1 U8551 ( .A(n8362), .Y(n8396) );
  INVX1 U8552 ( .A(n8362), .Y(n8397) );
  INVX1 U8553 ( .A(n8361), .Y(n8398) );
  INVX1 U8554 ( .A(n8361), .Y(n8399) );
  INVX1 U8555 ( .A(n8361), .Y(n8400) );
  INVX1 U8556 ( .A(n8360), .Y(n8401) );
  INVX1 U8557 ( .A(n8360), .Y(n8402) );
  INVX1 U8558 ( .A(n8360), .Y(n8403) );
  INVX1 U8559 ( .A(n8459), .Y(n8404) );
  INVX1 U8560 ( .A(n8370), .Y(n8405) );
  INVX1 U8561 ( .A(n8369), .Y(n8406) );
  INVX1 U8562 ( .A(n8359), .Y(n8407) );
  INVX1 U8563 ( .A(n8359), .Y(n8408) );
  INVX1 U8564 ( .A(n8359), .Y(n8409) );
  INVX1 U8565 ( .A(n8358), .Y(n8410) );
  INVX1 U8566 ( .A(n8358), .Y(n8411) );
  INVX1 U8567 ( .A(n8358), .Y(n8412) );
  INVX1 U8568 ( .A(n8357), .Y(n8413) );
  INVX1 U8569 ( .A(n8357), .Y(n8414) );
  INVX1 U8570 ( .A(n8357), .Y(n8415) );
  INVX1 U8571 ( .A(n8356), .Y(n8416) );
  INVX1 U8572 ( .A(n8356), .Y(n8417) );
  INVX1 U8573 ( .A(n8356), .Y(n8418) );
  INVX1 U8574 ( .A(n8355), .Y(n8419) );
  INVX1 U8575 ( .A(n8355), .Y(n8420) );
  INVX1 U8576 ( .A(n8355), .Y(n8421) );
  INVX1 U8577 ( .A(n8354), .Y(n8422) );
  INVX1 U8578 ( .A(n8354), .Y(n8423) );
  INVX1 U8579 ( .A(n8354), .Y(n8424) );
  INVX1 U8580 ( .A(n8356), .Y(n8425) );
  INVX1 U8581 ( .A(n8355), .Y(n8426) );
  INVX1 U8582 ( .A(n8354), .Y(n8427) );
  INVX1 U8583 ( .A(n8461), .Y(n8428) );
  INVX1 U8584 ( .A(n8358), .Y(n8429) );
  INVX1 U8585 ( .A(n8357), .Y(n8430) );
  INVX1 U8586 ( .A(n8364), .Y(n8431) );
  INVX1 U8587 ( .A(n8363), .Y(n8432) );
  INVX1 U8588 ( .A(n8362), .Y(n8433) );
  INVX1 U8589 ( .A(n10520), .Y(n10601) );
  INVX1 U8590 ( .A(n10520), .Y(n10602) );
  INVX1 U8591 ( .A(n10520), .Y(n10603) );
  INVX1 U8592 ( .A(n10520), .Y(n10604) );
  INVX1 U8593 ( .A(n10628), .Y(n10605) );
  INVX1 U8594 ( .A(n10526), .Y(n10606) );
  INVX1 U8595 ( .A(n10626), .Y(n10607) );
  INVX1 U8596 ( .A(n10624), .Y(n10608) );
  INVX1 U8597 ( .A(n10532), .Y(n10609) );
  INVX1 U8598 ( .A(n10519), .Y(n10610) );
  INVX1 U8599 ( .A(n10519), .Y(n10611) );
  INVX1 U8600 ( .A(n10519), .Y(n10612) );
  INVX1 U8601 ( .A(n10518), .Y(n10613) );
  INVX1 U8602 ( .A(n10518), .Y(n10614) );
  INVX1 U8603 ( .A(n10518), .Y(n10615) );
  INVX1 U8604 ( .A(n10627), .Y(n10616) );
  INVX1 U8605 ( .A(n10534), .Y(n10617) );
  INVX1 U8606 ( .A(n10533), .Y(n10618) );
  INVX1 U8607 ( .A(n8353), .Y(n8434) );
  INVX1 U8608 ( .A(n8353), .Y(n8435) );
  INVX1 U8609 ( .A(n8353), .Y(n8436) );
  INVX1 U8610 ( .A(n8353), .Y(n8437) );
  INVX1 U8611 ( .A(n8461), .Y(n8438) );
  INVX1 U8612 ( .A(n8359), .Y(n8439) );
  INVX1 U8613 ( .A(n8459), .Y(n8440) );
  INVX1 U8614 ( .A(n8457), .Y(n8441) );
  INVX1 U8615 ( .A(n8365), .Y(n8442) );
  INVX1 U8616 ( .A(n8352), .Y(n8443) );
  INVX1 U8617 ( .A(n8352), .Y(n8444) );
  INVX1 U8618 ( .A(n8352), .Y(n8445) );
  INVX1 U8619 ( .A(n8351), .Y(n8446) );
  INVX1 U8620 ( .A(n8351), .Y(n8447) );
  INVX1 U8621 ( .A(n8351), .Y(n8448) );
  INVX1 U8622 ( .A(n8460), .Y(n8449) );
  INVX1 U8623 ( .A(n8367), .Y(n8450) );
  INVX1 U8624 ( .A(n8366), .Y(n8451) );
  INVX1 U8625 ( .A(n10537), .Y(n10539) );
  INVX1 U8626 ( .A(n10537), .Y(n10540) );
  INVX1 U8627 ( .A(n10536), .Y(n10541) );
  INVX1 U8628 ( .A(n10536), .Y(n10542) );
  INVX1 U8629 ( .A(n10536), .Y(n10543) );
  INVX1 U8630 ( .A(n10535), .Y(n10544) );
  INVX1 U8631 ( .A(n10535), .Y(n10545) );
  INVX1 U8632 ( .A(n10535), .Y(n10546) );
  INVX1 U8633 ( .A(n8370), .Y(n8372) );
  INVX1 U8634 ( .A(n8370), .Y(n8373) );
  INVX1 U8635 ( .A(n8369), .Y(n8374) );
  INVX1 U8636 ( .A(n8369), .Y(n8375) );
  INVX1 U8637 ( .A(n8369), .Y(n8376) );
  INVX1 U8638 ( .A(n8368), .Y(n8377) );
  INVX1 U8639 ( .A(n8368), .Y(n8378) );
  INVX1 U8640 ( .A(n8368), .Y(n8379) );
  INVX1 U8641 ( .A(n10624), .Y(n10619) );
  INVX1 U8642 ( .A(n10519), .Y(n10620) );
  INVX1 U8643 ( .A(n10518), .Y(n10621) );
  INVX1 U8644 ( .A(n8457), .Y(n8452) );
  INVX1 U8645 ( .A(n8352), .Y(n8453) );
  INVX1 U8646 ( .A(n8351), .Y(n8454) );
  INVX1 U8647 ( .A(n10626), .Y(n10622) );
  INVX1 U8648 ( .A(n10624), .Y(n10623) );
  INVX1 U8649 ( .A(n8459), .Y(n8455) );
  INVX1 U8650 ( .A(n8457), .Y(n8456) );
  INVX1 U8651 ( .A(n10632), .Y(n10534) );
  INVX1 U8652 ( .A(n10632), .Y(n10533) );
  INVX1 U8653 ( .A(n10632), .Y(n10532) );
  INVX1 U8654 ( .A(n10631), .Y(n10531) );
  INVX1 U8655 ( .A(n10631), .Y(n10530) );
  INVX1 U8656 ( .A(n10631), .Y(n10529) );
  INVX1 U8657 ( .A(n10630), .Y(n10528) );
  INVX1 U8658 ( .A(n10629), .Y(n10527) );
  INVX1 U8659 ( .A(n10630), .Y(n10526) );
  INVX1 U8660 ( .A(n10630), .Y(n10525) );
  INVX1 U8661 ( .A(n10630), .Y(n10524) );
  INVX1 U8662 ( .A(n10629), .Y(n10523) );
  INVX1 U8663 ( .A(n10629), .Y(n10522) );
  INVX1 U8664 ( .A(n10629), .Y(n10521) );
  INVX1 U8665 ( .A(n8465), .Y(n8367) );
  INVX1 U8666 ( .A(n8465), .Y(n8366) );
  INVX1 U8667 ( .A(n8465), .Y(n8365) );
  INVX1 U8668 ( .A(n8464), .Y(n8364) );
  INVX1 U8669 ( .A(n8464), .Y(n8363) );
  INVX1 U8670 ( .A(n8464), .Y(n8362) );
  INVX1 U8671 ( .A(n8463), .Y(n8361) );
  INVX1 U8672 ( .A(n8462), .Y(n8360) );
  INVX1 U8673 ( .A(n8463), .Y(n8359) );
  INVX1 U8674 ( .A(n8463), .Y(n8358) );
  INVX1 U8675 ( .A(n8463), .Y(n8357) );
  INVX1 U8676 ( .A(n8462), .Y(n8356) );
  INVX1 U8677 ( .A(n8462), .Y(n8355) );
  INVX1 U8678 ( .A(n8462), .Y(n8354) );
  INVX1 U8679 ( .A(n10537), .Y(n10538) );
  INVX1 U8680 ( .A(n8370), .Y(n8371) );
  INVX1 U8681 ( .A(n10637), .Y(n10657) );
  INVX1 U8682 ( .A(n10682), .Y(n10658) );
  INVX1 U8683 ( .A(n10637), .Y(n10659) );
  INVX1 U8684 ( .A(n10634), .Y(n10660) );
  INVX1 U8685 ( .A(n10682), .Y(n10661) );
  INVX1 U8686 ( .A(n10635), .Y(n10662) );
  INVX1 U8687 ( .A(n10634), .Y(n10663) );
  INVX1 U8688 ( .A(n10635), .Y(n10664) );
  INVX1 U8689 ( .A(n10638), .Y(n10665) );
  INVX1 U8690 ( .A(n10634), .Y(n10666) );
  INVX1 U8691 ( .A(n10682), .Y(n10667) );
  INVX1 U8692 ( .A(n10635), .Y(n10668) );
  INVX1 U8693 ( .A(n10638), .Y(n10669) );
  INVX1 U8694 ( .A(n10682), .Y(n10670) );
  INVX1 U8695 ( .A(n10682), .Y(n10671) );
  INVX1 U8696 ( .A(n10682), .Y(n10672) );
  INVX1 U8697 ( .A(n10634), .Y(n10673) );
  INVX1 U8698 ( .A(n10636), .Y(n10674) );
  INVX1 U8699 ( .A(n10634), .Y(n10675) );
  INVX1 U8700 ( .A(n10638), .Y(n10676) );
  INVX1 U8701 ( .A(n10637), .Y(n10677) );
  INVX1 U8702 ( .A(n10682), .Y(n10678) );
  INVX1 U8703 ( .A(n10636), .Y(n10679) );
  INVX1 U8704 ( .A(n10636), .Y(n10680) );
  INVX1 U8705 ( .A(n8470), .Y(n8490) );
  INVX1 U8706 ( .A(n8515), .Y(n8491) );
  INVX1 U8707 ( .A(n8470), .Y(n8492) );
  INVX1 U8708 ( .A(n8467), .Y(n8493) );
  INVX1 U8709 ( .A(n8515), .Y(n8494) );
  INVX1 U8710 ( .A(n8468), .Y(n8495) );
  INVX1 U8711 ( .A(n8467), .Y(n8496) );
  INVX1 U8712 ( .A(n8468), .Y(n8497) );
  INVX1 U8713 ( .A(n8471), .Y(n8498) );
  INVX1 U8714 ( .A(n8467), .Y(n8499) );
  INVX1 U8715 ( .A(n8515), .Y(n8500) );
  INVX1 U8716 ( .A(n8468), .Y(n8501) );
  INVX1 U8717 ( .A(n8471), .Y(n8502) );
  INVX1 U8718 ( .A(n8515), .Y(n8503) );
  INVX1 U8719 ( .A(n8515), .Y(n8504) );
  INVX1 U8720 ( .A(n8515), .Y(n8505) );
  INVX1 U8721 ( .A(n8467), .Y(n8506) );
  INVX1 U8722 ( .A(n8469), .Y(n8507) );
  INVX1 U8723 ( .A(n8467), .Y(n8508) );
  INVX1 U8724 ( .A(n8471), .Y(n8509) );
  INVX1 U8725 ( .A(n8470), .Y(n8510) );
  INVX1 U8726 ( .A(n8515), .Y(n8511) );
  INVX1 U8727 ( .A(n8469), .Y(n8512) );
  INVX1 U8728 ( .A(n8469), .Y(n8513) );
  INVX1 U8729 ( .A(n10683), .Y(n10684) );
  INVX1 U8730 ( .A(n10683), .Y(n10685) );
  INVX1 U8731 ( .A(n10683), .Y(n10686) );
  INVX1 U8732 ( .A(n10683), .Y(n10687) );
  INVX1 U8733 ( .A(n10683), .Y(n10688) );
  INVX1 U8734 ( .A(n10683), .Y(n10689) );
  INVX1 U8735 ( .A(n10683), .Y(n10690) );
  INVX1 U8736 ( .A(n10683), .Y(n10691) );
  INVX1 U8737 ( .A(n10683), .Y(n10692) );
  INVX1 U8738 ( .A(n10683), .Y(n10693) );
  INVX1 U8739 ( .A(n10683), .Y(n10694) );
  INVX1 U8740 ( .A(n10683), .Y(n10695) );
  INVX1 U8741 ( .A(n10683), .Y(n10696) );
  INVX1 U8742 ( .A(n10683), .Y(n10697) );
  INVX1 U8743 ( .A(n10683), .Y(n10698) );
  INVX1 U8744 ( .A(n8516), .Y(n8517) );
  INVX1 U8745 ( .A(n8516), .Y(n8518) );
  INVX1 U8746 ( .A(n8516), .Y(n8519) );
  INVX1 U8747 ( .A(n8516), .Y(n8520) );
  INVX1 U8748 ( .A(n8516), .Y(n8521) );
  INVX1 U8749 ( .A(n8516), .Y(n8522) );
  INVX1 U8750 ( .A(n8516), .Y(n8523) );
  INVX1 U8751 ( .A(n8516), .Y(n8524) );
  INVX1 U8752 ( .A(n8516), .Y(n8525) );
  INVX1 U8753 ( .A(n8516), .Y(n8526) );
  INVX1 U8754 ( .A(n8516), .Y(n8527) );
  INVX1 U8755 ( .A(n8516), .Y(n8528) );
  INVX1 U8756 ( .A(n8516), .Y(n8529) );
  INVX1 U8757 ( .A(n8516), .Y(n8530) );
  INVX1 U8758 ( .A(n8516), .Y(n8531) );
  INVX1 U8759 ( .A(n10638), .Y(n10640) );
  INVX1 U8760 ( .A(n10638), .Y(n10641) );
  INVX1 U8761 ( .A(n10637), .Y(n10642) );
  INVX1 U8762 ( .A(n10637), .Y(n10643) );
  INVX1 U8763 ( .A(n10637), .Y(n10644) );
  INVX1 U8764 ( .A(n10635), .Y(n10645) );
  INVX1 U8765 ( .A(n10638), .Y(n10646) );
  INVX1 U8766 ( .A(n10637), .Y(n10647) );
  INVX1 U8767 ( .A(n10636), .Y(n10648) );
  INVX1 U8768 ( .A(n10636), .Y(n10649) );
  INVX1 U8769 ( .A(n10636), .Y(n10650) );
  INVX1 U8770 ( .A(n10635), .Y(n10651) );
  INVX1 U8771 ( .A(n10635), .Y(n10652) );
  INVX1 U8772 ( .A(n10635), .Y(n10653) );
  INVX1 U8773 ( .A(n10635), .Y(n10654) );
  INVX1 U8774 ( .A(n10634), .Y(n10655) );
  INVX1 U8775 ( .A(n10636), .Y(n10656) );
  INVX1 U8776 ( .A(n8471), .Y(n8473) );
  INVX1 U8777 ( .A(n8471), .Y(n8474) );
  INVX1 U8778 ( .A(n8470), .Y(n8475) );
  INVX1 U8779 ( .A(n8470), .Y(n8476) );
  INVX1 U8780 ( .A(n8470), .Y(n8477) );
  INVX1 U8781 ( .A(n8468), .Y(n8478) );
  INVX1 U8782 ( .A(n8471), .Y(n8479) );
  INVX1 U8783 ( .A(n8470), .Y(n8480) );
  INVX1 U8784 ( .A(n8469), .Y(n8481) );
  INVX1 U8785 ( .A(n8469), .Y(n8482) );
  INVX1 U8786 ( .A(n8469), .Y(n8483) );
  INVX1 U8787 ( .A(n8468), .Y(n8484) );
  INVX1 U8788 ( .A(n8468), .Y(n8485) );
  INVX1 U8789 ( .A(n8468), .Y(n8486) );
  INVX1 U8790 ( .A(n8468), .Y(n8487) );
  INVX1 U8791 ( .A(n8467), .Y(n8488) );
  INVX1 U8792 ( .A(n8469), .Y(n8489) );
  INVX1 U8793 ( .A(n10683), .Y(n10699) );
  INVX1 U8794 ( .A(n10683), .Y(n10700) );
  INVX1 U8795 ( .A(n8516), .Y(n8532) );
  INVX1 U8796 ( .A(n8516), .Y(n8533) );
  INVX1 U8797 ( .A(n166), .Y(n10764) );
  INVX1 U8798 ( .A(n233), .Y(n10762) );
  INVX1 U8799 ( .A(n299), .Y(n10760) );
  INVX1 U8800 ( .A(n365), .Y(n10758) );
  INVX1 U8801 ( .A(n431), .Y(n10756) );
  INVX1 U8802 ( .A(n497), .Y(n10754) );
  INVX1 U8803 ( .A(n563), .Y(n10752) );
  INVX1 U8804 ( .A(n696), .Y(n10748) );
  INVX1 U8805 ( .A(n762), .Y(n10746) );
  INVX1 U8806 ( .A(n827), .Y(n10744) );
  INVX1 U8807 ( .A(n892), .Y(n10742) );
  INVX1 U8808 ( .A(n957), .Y(n10740) );
  INVX1 U8809 ( .A(n1022), .Y(n10738) );
  INVX1 U8810 ( .A(n1087), .Y(n10736) );
  INVX1 U8811 ( .A(n1283), .Y(n10730) );
  INVX1 U8812 ( .A(n1738), .Y(n10716) );
  INVX1 U8813 ( .A(n1478), .Y(n10724) );
  INVX1 U8814 ( .A(n1543), .Y(n10722) );
  INVX1 U8815 ( .A(n1608), .Y(n10720) );
  INVX1 U8816 ( .A(n1673), .Y(n10718) );
  INVX1 U8817 ( .A(n1804), .Y(n10714) );
  INVX1 U8818 ( .A(n1869), .Y(n10712) );
  INVX1 U8819 ( .A(n2064), .Y(n10706) );
  INVX1 U8820 ( .A(n10638), .Y(n10639) );
  INVX1 U8821 ( .A(n8471), .Y(n8472) );
  INVX1 U8822 ( .A(n10627), .Y(n10632) );
  INVX1 U8823 ( .A(n10627), .Y(n10631) );
  INVX1 U8824 ( .A(n10628), .Y(n10630) );
  INVX1 U8825 ( .A(n10628), .Y(n10629) );
  INVX1 U8826 ( .A(n8460), .Y(n8465) );
  INVX1 U8827 ( .A(n8460), .Y(n8464) );
  INVX1 U8828 ( .A(n8461), .Y(n8463) );
  INVX1 U8829 ( .A(n8461), .Y(n8462) );
  INVX1 U8830 ( .A(n10625), .Y(n10520) );
  INVX1 U8831 ( .A(N18), .Y(n10519) );
  INVX1 U8832 ( .A(N18), .Y(n10518) );
  INVX1 U8833 ( .A(n8458), .Y(n8353) );
  INVX1 U8834 ( .A(N13), .Y(n8352) );
  INVX1 U8835 ( .A(N13), .Y(n8351) );
  INVX1 U8836 ( .A(n10633), .Y(n10537) );
  INVX1 U8837 ( .A(n10633), .Y(n10536) );
  INVX1 U8838 ( .A(n10633), .Y(n10535) );
  INVX1 U8839 ( .A(n8466), .Y(n8370) );
  INVX1 U8840 ( .A(n8466), .Y(n8369) );
  INVX1 U8841 ( .A(n8466), .Y(n8368) );
  INVX1 U8842 ( .A(n10766), .Y(n10765) );
  INVX1 U8843 ( .A(n10634), .Y(n10681) );
  INVX1 U8844 ( .A(N19), .Y(n10634) );
  INVX1 U8845 ( .A(n8467), .Y(n8514) );
  INVX1 U8846 ( .A(N14), .Y(n8467) );
  INVX1 U8847 ( .A(n629), .Y(n10750) );
  INVX1 U8848 ( .A(n1152), .Y(n10734) );
  INVX1 U8849 ( .A(n1217), .Y(n10732) );
  INVX1 U8850 ( .A(n1348), .Y(n10728) );
  INVX1 U8851 ( .A(n1413), .Y(n10726) );
  INVX1 U8852 ( .A(n1934), .Y(n10710) );
  INVX1 U8853 ( .A(n1999), .Y(n10708) );
  INVX1 U8854 ( .A(n2129), .Y(n10704) );
  INVX1 U8855 ( .A(n2194), .Y(n10702) );
  INVX1 U8856 ( .A(N20), .Y(n10683) );
  INVX1 U8857 ( .A(N15), .Y(n8516) );
  INVX1 U8858 ( .A(n166), .Y(n10763) );
  INVX1 U8859 ( .A(n233), .Y(n10761) );
  INVX1 U8860 ( .A(n299), .Y(n10759) );
  INVX1 U8861 ( .A(n365), .Y(n10757) );
  INVX1 U8862 ( .A(n431), .Y(n10755) );
  INVX1 U8863 ( .A(n497), .Y(n10753) );
  INVX1 U8864 ( .A(n563), .Y(n10751) );
  INVX1 U8865 ( .A(n629), .Y(n10749) );
  INVX1 U8866 ( .A(n696), .Y(n10747) );
  INVX1 U8867 ( .A(n1217), .Y(n10731) );
  INVX1 U8868 ( .A(n1738), .Y(n10715) );
  INVX1 U8869 ( .A(n762), .Y(n10745) );
  INVX1 U8870 ( .A(n827), .Y(n10743) );
  INVX1 U8871 ( .A(n892), .Y(n10741) );
  INVX1 U8872 ( .A(n957), .Y(n10739) );
  INVX1 U8873 ( .A(n1022), .Y(n10737) );
  INVX1 U8874 ( .A(n1087), .Y(n10735) );
  INVX1 U8875 ( .A(n1152), .Y(n10733) );
  INVX1 U8876 ( .A(n1283), .Y(n10729) );
  INVX1 U8877 ( .A(n1348), .Y(n10727) );
  INVX1 U8878 ( .A(n1413), .Y(n10725) );
  INVX1 U8879 ( .A(n1478), .Y(n10723) );
  INVX1 U8880 ( .A(n1543), .Y(n10721) );
  INVX1 U8881 ( .A(n1608), .Y(n10719) );
  INVX1 U8882 ( .A(n1673), .Y(n10717) );
  INVX1 U8883 ( .A(n1804), .Y(n10713) );
  INVX1 U8884 ( .A(n1869), .Y(n10711) );
  INVX1 U8885 ( .A(n1934), .Y(n10709) );
  INVX1 U8886 ( .A(n1999), .Y(n10707) );
  INVX1 U8887 ( .A(n2064), .Y(n10705) );
  INVX1 U8888 ( .A(n2129), .Y(n10703) );
  INVX1 U8889 ( .A(n2194), .Y(n10701) );
  INVX1 U8890 ( .A(n10625), .Y(n10627) );
  INVX1 U8891 ( .A(n10625), .Y(n10628) );
  INVX1 U8892 ( .A(n8458), .Y(n8460) );
  INVX1 U8893 ( .A(n8458), .Y(n8461) );
  INVX1 U8894 ( .A(N19), .Y(n10638) );
  INVX1 U8895 ( .A(N19), .Y(n10637) );
  INVX1 U8896 ( .A(N19), .Y(n10636) );
  INVX1 U8897 ( .A(N19), .Y(n10635) );
  INVX1 U8898 ( .A(N14), .Y(n8471) );
  INVX1 U8899 ( .A(N14), .Y(n8470) );
  INVX1 U8900 ( .A(N14), .Y(n8469) );
  INVX1 U8901 ( .A(N14), .Y(n8468) );
  INVX1 U8902 ( .A(n10626), .Y(n10633) );
  INVX1 U8903 ( .A(n10625), .Y(n10626) );
  INVX1 U8904 ( .A(n8459), .Y(n8466) );
  INVX1 U8905 ( .A(n8458), .Y(n8459) );
  INVX1 U8906 ( .A(n6303), .Y(n10830) );
  INVX1 U8907 ( .A(n6304), .Y(n10779) );
  INVX1 U8908 ( .A(n6305), .Y(n10778) );
  INVX1 U8909 ( .A(n6306), .Y(n10777) );
  INVX1 U8910 ( .A(n6307), .Y(n10776) );
  INVX1 U8911 ( .A(n6308), .Y(n10775) );
  INVX1 U8912 ( .A(n6309), .Y(n10774) );
  INVX1 U8913 ( .A(n6310), .Y(n10773) );
  INVX1 U8914 ( .A(n6311), .Y(n10772) );
  INVX1 U8915 ( .A(n6312), .Y(n10771) );
  INVX1 U8916 ( .A(n6313), .Y(n10770) );
  INVX1 U8917 ( .A(n6314), .Y(n10769) );
  INVX1 U8918 ( .A(n6315), .Y(n10768) );
  INVX1 U8919 ( .A(n6316), .Y(n10829) );
  INVX1 U8920 ( .A(n6317), .Y(n10828) );
  INVX1 U8921 ( .A(n6318), .Y(n10827) );
  INVX1 U8922 ( .A(n6319), .Y(n10826) );
  INVX1 U8923 ( .A(n6320), .Y(n10825) );
  INVX1 U8924 ( .A(n6321), .Y(n10824) );
  INVX1 U8925 ( .A(n6322), .Y(n10823) );
  INVX1 U8926 ( .A(n6323), .Y(n10822) );
  INVX1 U8927 ( .A(n6324), .Y(n10821) );
  INVX1 U8928 ( .A(n6325), .Y(n10820) );
  INVX1 U8929 ( .A(n6326), .Y(n10819) );
  INVX1 U8930 ( .A(n6327), .Y(n10818) );
  INVX1 U8931 ( .A(n6328), .Y(n10817) );
  INVX1 U8932 ( .A(n6329), .Y(n10816) );
  INVX1 U8933 ( .A(n6330), .Y(n10815) );
  INVX1 U8934 ( .A(n6331), .Y(n10814) );
  INVX1 U8935 ( .A(n6332), .Y(n10813) );
  INVX1 U8936 ( .A(n6333), .Y(n10812) );
  INVX1 U8937 ( .A(n6334), .Y(n10811) );
  INVX1 U8938 ( .A(n6335), .Y(n10810) );
  INVX1 U8939 ( .A(n6336), .Y(n10809) );
  INVX1 U8940 ( .A(n6337), .Y(n10808) );
  INVX1 U8941 ( .A(n6338), .Y(n10807) );
  INVX1 U8942 ( .A(n6339), .Y(n10806) );
  INVX1 U8943 ( .A(n6340), .Y(n10805) );
  INVX1 U8944 ( .A(n6341), .Y(n10804) );
  INVX1 U8945 ( .A(n6342), .Y(n10803) );
  INVX1 U8946 ( .A(n6343), .Y(n10802) );
  INVX1 U8947 ( .A(n6344), .Y(n10801) );
  INVX1 U8948 ( .A(n6345), .Y(n10800) );
  INVX1 U8949 ( .A(n6346), .Y(n10799) );
  INVX1 U8950 ( .A(n6347), .Y(n10798) );
  INVX1 U8951 ( .A(n6348), .Y(n10797) );
  INVX1 U8952 ( .A(n6349), .Y(n10796) );
  INVX1 U8953 ( .A(n6350), .Y(n10795) );
  INVX1 U8954 ( .A(n6351), .Y(n10794) );
  INVX1 U8955 ( .A(n6352), .Y(n10793) );
  INVX1 U8956 ( .A(n6353), .Y(n10792) );
  INVX1 U8957 ( .A(n6354), .Y(n10791) );
  INVX1 U8958 ( .A(n6355), .Y(n10790) );
  INVX1 U8959 ( .A(n6356), .Y(n10789) );
  INVX1 U8960 ( .A(n6357), .Y(n10788) );
  INVX1 U8961 ( .A(n6358), .Y(n10787) );
  INVX1 U8962 ( .A(n6359), .Y(n10786) );
  INVX1 U8963 ( .A(n6360), .Y(n10785) );
  INVX1 U8964 ( .A(n6361), .Y(n10784) );
  INVX1 U8965 ( .A(n6362), .Y(n10783) );
  INVX1 U8966 ( .A(n6363), .Y(n10782) );
  INVX1 U8967 ( .A(n6364), .Y(n10781) );
  INVX1 U8968 ( .A(n6365), .Y(n10780) );
  INVX1 U8969 ( .A(n6366), .Y(n10767) );
  INVX1 U8970 ( .A(n631), .Y(n10766) );
  INVX1 U8971 ( .A(n10624), .Y(n10625) );
  INVX1 U8972 ( .A(n8457), .Y(n8458) );
  AND2X1 U8973 ( .A(write_en), .B(reset_n), .Y(n631) );
  AND2X1 U8974 ( .A(wdata[0]), .B(n631), .Y(n6303) );
  AND2X1 U8975 ( .A(wdata[51]), .B(n10765), .Y(n6304) );
  AND2X1 U8976 ( .A(wdata[52]), .B(n631), .Y(n6305) );
  AND2X1 U8977 ( .A(wdata[53]), .B(n631), .Y(n6306) );
  AND2X1 U8978 ( .A(wdata[54]), .B(n10765), .Y(n6307) );
  AND2X1 U8979 ( .A(wdata[55]), .B(n631), .Y(n6308) );
  AND2X1 U8980 ( .A(wdata[56]), .B(n631), .Y(n6309) );
  AND2X1 U8981 ( .A(wdata[57]), .B(n10765), .Y(n6310) );
  AND2X1 U8982 ( .A(wdata[58]), .B(n10765), .Y(n6311) );
  AND2X1 U8983 ( .A(wdata[59]), .B(n631), .Y(n6312) );
  AND2X1 U8984 ( .A(wdata[60]), .B(n10765), .Y(n6313) );
  AND2X1 U8985 ( .A(wdata[61]), .B(n631), .Y(n6314) );
  AND2X1 U8986 ( .A(wdata[62]), .B(n631), .Y(n6315) );
  AND2X1 U8987 ( .A(wdata[1]), .B(n631), .Y(n6316) );
  AND2X1 U8988 ( .A(wdata[2]), .B(n631), .Y(n6317) );
  AND2X1 U8989 ( .A(wdata[3]), .B(n631), .Y(n6318) );
  AND2X1 U8990 ( .A(wdata[4]), .B(n631), .Y(n6319) );
  AND2X1 U8991 ( .A(wdata[5]), .B(n631), .Y(n6320) );
  AND2X1 U8992 ( .A(wdata[6]), .B(n631), .Y(n6321) );
  AND2X1 U8993 ( .A(wdata[7]), .B(n631), .Y(n6322) );
  AND2X1 U8994 ( .A(wdata[8]), .B(n631), .Y(n6323) );
  AND2X1 U8995 ( .A(wdata[9]), .B(n631), .Y(n6324) );
  AND2X1 U8996 ( .A(wdata[10]), .B(n631), .Y(n6325) );
  AND2X1 U8997 ( .A(wdata[11]), .B(n631), .Y(n6326) );
  AND2X1 U8998 ( .A(wdata[12]), .B(n631), .Y(n6327) );
  AND2X1 U8999 ( .A(wdata[13]), .B(n631), .Y(n6328) );
  AND2X1 U9000 ( .A(wdata[14]), .B(n631), .Y(n6329) );
  AND2X1 U9001 ( .A(wdata[15]), .B(n631), .Y(n6330) );
  AND2X1 U9002 ( .A(wdata[16]), .B(n10765), .Y(n6331) );
  AND2X1 U9003 ( .A(wdata[17]), .B(n10765), .Y(n6332) );
  AND2X1 U9004 ( .A(wdata[18]), .B(n10765), .Y(n6333) );
  AND2X1 U9005 ( .A(wdata[19]), .B(n10765), .Y(n6334) );
  AND2X1 U9006 ( .A(wdata[20]), .B(n10765), .Y(n6335) );
  AND2X1 U9007 ( .A(wdata[21]), .B(n10765), .Y(n6336) );
  AND2X1 U9008 ( .A(wdata[22]), .B(n10765), .Y(n6337) );
  AND2X1 U9009 ( .A(wdata[23]), .B(n10765), .Y(n6338) );
  AND2X1 U9010 ( .A(wdata[24]), .B(n10765), .Y(n6339) );
  AND2X1 U9011 ( .A(wdata[25]), .B(n10765), .Y(n6340) );
  AND2X1 U9012 ( .A(wdata[26]), .B(n10765), .Y(n6341) );
  AND2X1 U9013 ( .A(wdata[27]), .B(n10765), .Y(n6342) );
  AND2X1 U9014 ( .A(wdata[28]), .B(n10765), .Y(n6343) );
  AND2X1 U9015 ( .A(wdata[29]), .B(n10765), .Y(n6344) );
  AND2X1 U9016 ( .A(wdata[30]), .B(n10765), .Y(n6345) );
  AND2X1 U9017 ( .A(wdata[31]), .B(n10765), .Y(n6346) );
  AND2X1 U9018 ( .A(wdata[32]), .B(n10765), .Y(n6347) );
  AND2X1 U9019 ( .A(wdata[33]), .B(n10765), .Y(n6348) );
  AND2X1 U9020 ( .A(wdata[34]), .B(n631), .Y(n6349) );
  AND2X1 U9021 ( .A(wdata[35]), .B(n10765), .Y(n6350) );
  AND2X1 U9022 ( .A(wdata[36]), .B(n631), .Y(n6351) );
  AND2X1 U9023 ( .A(wdata[37]), .B(n10765), .Y(n6352) );
  AND2X1 U9024 ( .A(wdata[38]), .B(n631), .Y(n6353) );
  AND2X1 U9025 ( .A(wdata[39]), .B(n10765), .Y(n6354) );
  AND2X1 U9026 ( .A(wdata[40]), .B(n631), .Y(n6355) );
  AND2X1 U9027 ( .A(wdata[41]), .B(n10765), .Y(n6356) );
  AND2X1 U9028 ( .A(wdata[42]), .B(n631), .Y(n6357) );
  AND2X1 U9029 ( .A(wdata[43]), .B(n10765), .Y(n6358) );
  AND2X1 U9030 ( .A(wdata[44]), .B(n631), .Y(n6359) );
  AND2X1 U9031 ( .A(wdata[45]), .B(n10765), .Y(n6360) );
  AND2X1 U9032 ( .A(wdata[46]), .B(n631), .Y(n6361) );
  AND2X1 U9033 ( .A(wdata[47]), .B(n10765), .Y(n6362) );
  AND2X1 U9034 ( .A(wdata[48]), .B(n10765), .Y(n6363) );
  AND2X1 U9035 ( .A(wdata[49]), .B(n631), .Y(n6364) );
  AND2X1 U9036 ( .A(wdata[50]), .B(n10765), .Y(n6365) );
  AND2X1 U9037 ( .A(wdata[63]), .B(n631), .Y(n6366) );
  INVX1 U9038 ( .A(waddr[2]), .Y(n10833) );
  INVX1 U9039 ( .A(waddr[0]), .Y(n10835) );
  INVX1 U9040 ( .A(waddr[1]), .Y(n10834) );
  INVX1 U9041 ( .A(N19), .Y(n10682) );
  INVX1 U9042 ( .A(N14), .Y(n8515) );
  INVX1 U9043 ( .A(N18), .Y(n10624) );
  INVX1 U9044 ( .A(N13), .Y(n8457) );
  AND2X1 U9045 ( .A(N152), .B(read_en[1]), .Y(rdata_1[0]) );
  INVX1 U9046 ( .A(n10454), .Y(N152) );
  AND2X1 U9047 ( .A(N151), .B(read_en[1]), .Y(rdata_1[1]) );
  INVX1 U9048 ( .A(n10455), .Y(N151) );
  AND2X1 U9049 ( .A(N150), .B(read_en[1]), .Y(rdata_1[2]) );
  INVX1 U9050 ( .A(n10456), .Y(N150) );
  AND2X1 U9051 ( .A(N149), .B(read_en[1]), .Y(rdata_1[3]) );
  INVX1 U9052 ( .A(n10457), .Y(N149) );
  AND2X1 U9053 ( .A(N148), .B(read_en[1]), .Y(rdata_1[4]) );
  INVX1 U9054 ( .A(n10458), .Y(N148) );
  AND2X1 U9055 ( .A(N147), .B(read_en[1]), .Y(rdata_1[5]) );
  INVX1 U9056 ( .A(n10459), .Y(N147) );
  AND2X1 U9057 ( .A(N146), .B(read_en[1]), .Y(rdata_1[6]) );
  INVX1 U9058 ( .A(n10460), .Y(N146) );
  AND2X1 U9059 ( .A(N145), .B(read_en[1]), .Y(rdata_1[7]) );
  INVX1 U9060 ( .A(n10461), .Y(N145) );
  AND2X1 U9061 ( .A(N144), .B(read_en[1]), .Y(rdata_1[8]) );
  INVX1 U9062 ( .A(n10462), .Y(N144) );
  AND2X1 U9063 ( .A(read_en[1]), .B(N143), .Y(rdata_1[9]) );
  INVX1 U9064 ( .A(n10463), .Y(N143) );
  AND2X1 U9065 ( .A(N142), .B(read_en[1]), .Y(rdata_1[10]) );
  INVX1 U9066 ( .A(n10464), .Y(N142) );
  AND2X1 U9067 ( .A(N141), .B(read_en[1]), .Y(rdata_1[11]) );
  INVX1 U9068 ( .A(n10465), .Y(N141) );
  AND2X1 U9069 ( .A(N140), .B(read_en[1]), .Y(rdata_1[12]) );
  INVX1 U9070 ( .A(n10466), .Y(N140) );
  AND2X1 U9071 ( .A(N139), .B(read_en[1]), .Y(rdata_1[13]) );
  INVX1 U9072 ( .A(n10467), .Y(N139) );
  AND2X1 U9073 ( .A(N138), .B(read_en[1]), .Y(rdata_1[14]) );
  INVX1 U9074 ( .A(n10468), .Y(N138) );
  AND2X1 U9075 ( .A(N137), .B(read_en[1]), .Y(rdata_1[15]) );
  INVX1 U9076 ( .A(n10469), .Y(N137) );
  AND2X1 U9077 ( .A(N136), .B(read_en[1]), .Y(rdata_1[16]) );
  INVX1 U9078 ( .A(n10470), .Y(N136) );
  AND2X1 U9079 ( .A(N135), .B(read_en[1]), .Y(rdata_1[17]) );
  INVX1 U9080 ( .A(n10471), .Y(N135) );
  AND2X1 U9081 ( .A(N134), .B(read_en[1]), .Y(rdata_1[18]) );
  INVX1 U9082 ( .A(n10472), .Y(N134) );
  AND2X1 U9083 ( .A(N133), .B(read_en[1]), .Y(rdata_1[19]) );
  INVX1 U9084 ( .A(n10473), .Y(N133) );
  AND2X1 U9085 ( .A(N132), .B(read_en[1]), .Y(rdata_1[20]) );
  INVX1 U9086 ( .A(n10474), .Y(N132) );
  AND2X1 U9087 ( .A(N131), .B(read_en[1]), .Y(rdata_1[21]) );
  INVX1 U9088 ( .A(n10475), .Y(N131) );
  AND2X1 U9089 ( .A(N130), .B(read_en[1]), .Y(rdata_1[22]) );
  INVX1 U9090 ( .A(n10476), .Y(N130) );
  AND2X1 U9091 ( .A(N129), .B(read_en[1]), .Y(rdata_1[23]) );
  INVX1 U9092 ( .A(n10477), .Y(N129) );
  AND2X1 U9093 ( .A(N128), .B(read_en[1]), .Y(rdata_1[24]) );
  INVX1 U9094 ( .A(n10478), .Y(N128) );
  AND2X1 U9095 ( .A(N127), .B(read_en[1]), .Y(rdata_1[25]) );
  INVX1 U9096 ( .A(n10479), .Y(N127) );
  AND2X1 U9097 ( .A(N126), .B(read_en[1]), .Y(rdata_1[26]) );
  INVX1 U9098 ( .A(n10480), .Y(N126) );
  AND2X1 U9099 ( .A(N125), .B(read_en[1]), .Y(rdata_1[27]) );
  INVX1 U9100 ( .A(n10481), .Y(N125) );
  AND2X1 U9101 ( .A(N124), .B(read_en[1]), .Y(rdata_1[28]) );
  INVX1 U9102 ( .A(n10482), .Y(N124) );
  AND2X1 U9103 ( .A(N123), .B(read_en[1]), .Y(rdata_1[29]) );
  INVX1 U9104 ( .A(n10483), .Y(N123) );
  AND2X1 U9105 ( .A(N122), .B(read_en[1]), .Y(rdata_1[30]) );
  INVX1 U9106 ( .A(n10484), .Y(N122) );
  AND2X1 U9107 ( .A(N121), .B(read_en[1]), .Y(rdata_1[31]) );
  INVX1 U9108 ( .A(n10485), .Y(N121) );
  AND2X1 U9109 ( .A(N120), .B(read_en[1]), .Y(rdata_1[32]) );
  INVX1 U9110 ( .A(n10486), .Y(N120) );
  AND2X1 U9111 ( .A(N119), .B(read_en[1]), .Y(rdata_1[33]) );
  INVX1 U9112 ( .A(n10487), .Y(N119) );
  AND2X1 U9113 ( .A(N118), .B(read_en[1]), .Y(rdata_1[34]) );
  INVX1 U9114 ( .A(n10488), .Y(N118) );
  AND2X1 U9115 ( .A(N117), .B(read_en[1]), .Y(rdata_1[35]) );
  INVX1 U9116 ( .A(n10489), .Y(N117) );
  AND2X1 U9117 ( .A(N116), .B(read_en[1]), .Y(rdata_1[36]) );
  INVX1 U9118 ( .A(n10490), .Y(N116) );
  AND2X1 U9119 ( .A(N115), .B(read_en[1]), .Y(rdata_1[37]) );
  INVX1 U9120 ( .A(n10491), .Y(N115) );
  AND2X1 U9121 ( .A(N114), .B(read_en[1]), .Y(rdata_1[38]) );
  INVX1 U9122 ( .A(n10492), .Y(N114) );
  AND2X1 U9123 ( .A(N113), .B(read_en[1]), .Y(rdata_1[39]) );
  INVX1 U9124 ( .A(n10493), .Y(N113) );
  AND2X1 U9125 ( .A(N112), .B(read_en[1]), .Y(rdata_1[40]) );
  INVX1 U9126 ( .A(n10494), .Y(N112) );
  AND2X1 U9127 ( .A(N111), .B(read_en[1]), .Y(rdata_1[41]) );
  INVX1 U9128 ( .A(n10495), .Y(N111) );
  AND2X1 U9129 ( .A(N110), .B(read_en[1]), .Y(rdata_1[42]) );
  INVX1 U9130 ( .A(n10496), .Y(N110) );
  AND2X1 U9131 ( .A(N109), .B(read_en[1]), .Y(rdata_1[43]) );
  INVX1 U9132 ( .A(n10497), .Y(N109) );
  AND2X1 U9133 ( .A(N108), .B(read_en[1]), .Y(rdata_1[44]) );
  INVX1 U9134 ( .A(n10498), .Y(N108) );
  AND2X1 U9135 ( .A(N107), .B(read_en[1]), .Y(rdata_1[45]) );
  INVX1 U9136 ( .A(n10499), .Y(N107) );
  AND2X1 U9137 ( .A(N106), .B(read_en[1]), .Y(rdata_1[46]) );
  INVX1 U9138 ( .A(n10500), .Y(N106) );
  AND2X1 U9139 ( .A(N105), .B(read_en[1]), .Y(rdata_1[47]) );
  INVX1 U9140 ( .A(n10501), .Y(N105) );
  AND2X1 U9141 ( .A(N104), .B(read_en[1]), .Y(rdata_1[48]) );
  INVX1 U9142 ( .A(n10502), .Y(N104) );
  AND2X1 U9143 ( .A(N103), .B(read_en[1]), .Y(rdata_1[49]) );
  INVX1 U9144 ( .A(n10503), .Y(N103) );
  AND2X1 U9145 ( .A(N102), .B(read_en[1]), .Y(rdata_1[50]) );
  INVX1 U9146 ( .A(n10504), .Y(N102) );
  AND2X1 U9147 ( .A(N101), .B(read_en[1]), .Y(rdata_1[51]) );
  INVX1 U9148 ( .A(n10505), .Y(N101) );
  AND2X1 U9149 ( .A(N100), .B(read_en[1]), .Y(rdata_1[52]) );
  INVX1 U9150 ( .A(n10506), .Y(N100) );
  AND2X1 U9151 ( .A(N99), .B(read_en[1]), .Y(rdata_1[53]) );
  INVX1 U9152 ( .A(n10507), .Y(N99) );
  AND2X1 U9153 ( .A(N98), .B(read_en[1]), .Y(rdata_1[54]) );
  INVX1 U9154 ( .A(n10508), .Y(N98) );
  AND2X1 U9155 ( .A(N97), .B(read_en[1]), .Y(rdata_1[55]) );
  INVX1 U9156 ( .A(n10509), .Y(N97) );
  AND2X1 U9157 ( .A(N96), .B(read_en[1]), .Y(rdata_1[56]) );
  INVX1 U9158 ( .A(n10510), .Y(N96) );
  AND2X1 U9159 ( .A(N95), .B(read_en[1]), .Y(rdata_1[57]) );
  INVX1 U9160 ( .A(n10511), .Y(N95) );
  AND2X1 U9161 ( .A(N94), .B(read_en[1]), .Y(rdata_1[58]) );
  INVX1 U9162 ( .A(n10512), .Y(N94) );
  AND2X1 U9163 ( .A(N93), .B(read_en[1]), .Y(rdata_1[59]) );
  INVX1 U9164 ( .A(n10513), .Y(N93) );
  AND2X1 U9165 ( .A(N92), .B(read_en[1]), .Y(rdata_1[60]) );
  INVX1 U9166 ( .A(n10514), .Y(N92) );
  AND2X1 U9167 ( .A(N91), .B(read_en[1]), .Y(rdata_1[61]) );
  INVX1 U9168 ( .A(n10515), .Y(N91) );
  AND2X1 U9169 ( .A(N90), .B(read_en[1]), .Y(rdata_1[62]) );
  INVX1 U9170 ( .A(n10516), .Y(N90) );
  AND2X1 U9171 ( .A(N89), .B(read_en[1]), .Y(rdata_1[63]) );
  INVX1 U9172 ( .A(n10517), .Y(N89) );
  AND2X1 U9173 ( .A(N87), .B(read_en[0]), .Y(rdata_0[0]) );
  INVX1 U9174 ( .A(n8287), .Y(N87) );
  AND2X1 U9175 ( .A(N86), .B(read_en[0]), .Y(rdata_0[1]) );
  INVX1 U9176 ( .A(n8288), .Y(N86) );
  AND2X1 U9177 ( .A(N85), .B(read_en[0]), .Y(rdata_0[2]) );
  INVX1 U9178 ( .A(n8289), .Y(N85) );
  AND2X1 U9179 ( .A(N84), .B(read_en[0]), .Y(rdata_0[3]) );
  INVX1 U9180 ( .A(n8290), .Y(N84) );
  AND2X1 U9181 ( .A(N83), .B(read_en[0]), .Y(rdata_0[4]) );
  INVX1 U9182 ( .A(n8291), .Y(N83) );
  AND2X1 U9183 ( .A(N82), .B(read_en[0]), .Y(rdata_0[5]) );
  INVX1 U9184 ( .A(n8292), .Y(N82) );
  AND2X1 U9185 ( .A(N81), .B(read_en[0]), .Y(rdata_0[6]) );
  INVX1 U9186 ( .A(n8293), .Y(N81) );
  AND2X1 U9187 ( .A(N80), .B(read_en[0]), .Y(rdata_0[7]) );
  INVX1 U9188 ( .A(n8294), .Y(N80) );
  AND2X1 U9189 ( .A(N79), .B(read_en[0]), .Y(rdata_0[8]) );
  INVX1 U9190 ( .A(n8295), .Y(N79) );
  AND2X1 U9191 ( .A(read_en[0]), .B(N78), .Y(rdata_0[9]) );
  INVX1 U9192 ( .A(n8296), .Y(N78) );
  AND2X1 U9193 ( .A(N77), .B(read_en[0]), .Y(rdata_0[10]) );
  INVX1 U9194 ( .A(n8297), .Y(N77) );
  AND2X1 U9195 ( .A(N76), .B(read_en[0]), .Y(rdata_0[11]) );
  INVX1 U9196 ( .A(n8298), .Y(N76) );
  AND2X1 U9197 ( .A(N75), .B(read_en[0]), .Y(rdata_0[12]) );
  INVX1 U9198 ( .A(n8299), .Y(N75) );
  AND2X1 U9199 ( .A(N74), .B(read_en[0]), .Y(rdata_0[13]) );
  INVX1 U9200 ( .A(n8300), .Y(N74) );
  AND2X1 U9201 ( .A(N73), .B(read_en[0]), .Y(rdata_0[14]) );
  INVX1 U9202 ( .A(n8301), .Y(N73) );
  AND2X1 U9203 ( .A(N72), .B(read_en[0]), .Y(rdata_0[15]) );
  INVX1 U9204 ( .A(n8302), .Y(N72) );
  AND2X1 U9205 ( .A(N71), .B(read_en[0]), .Y(rdata_0[16]) );
  INVX1 U9206 ( .A(n8303), .Y(N71) );
  AND2X1 U9207 ( .A(N70), .B(read_en[0]), .Y(rdata_0[17]) );
  INVX1 U9208 ( .A(n8304), .Y(N70) );
  AND2X1 U9209 ( .A(N69), .B(read_en[0]), .Y(rdata_0[18]) );
  INVX1 U9210 ( .A(n8305), .Y(N69) );
  AND2X1 U9211 ( .A(N68), .B(read_en[0]), .Y(rdata_0[19]) );
  INVX1 U9212 ( .A(n8306), .Y(N68) );
  AND2X1 U9213 ( .A(N67), .B(read_en[0]), .Y(rdata_0[20]) );
  INVX1 U9214 ( .A(n8307), .Y(N67) );
  AND2X1 U9215 ( .A(N66), .B(read_en[0]), .Y(rdata_0[21]) );
  INVX1 U9216 ( .A(n8308), .Y(N66) );
  AND2X1 U9217 ( .A(N65), .B(read_en[0]), .Y(rdata_0[22]) );
  INVX1 U9218 ( .A(n8309), .Y(N65) );
  AND2X1 U9219 ( .A(N64), .B(read_en[0]), .Y(rdata_0[23]) );
  INVX1 U9220 ( .A(n8310), .Y(N64) );
  AND2X1 U9221 ( .A(N63), .B(read_en[0]), .Y(rdata_0[24]) );
  INVX1 U9222 ( .A(n8311), .Y(N63) );
  AND2X1 U9223 ( .A(N62), .B(read_en[0]), .Y(rdata_0[25]) );
  INVX1 U9224 ( .A(n8312), .Y(N62) );
  AND2X1 U9225 ( .A(N61), .B(read_en[0]), .Y(rdata_0[26]) );
  INVX1 U9226 ( .A(n8313), .Y(N61) );
  AND2X1 U9227 ( .A(N60), .B(read_en[0]), .Y(rdata_0[27]) );
  INVX1 U9228 ( .A(n8314), .Y(N60) );
  AND2X1 U9229 ( .A(N59), .B(read_en[0]), .Y(rdata_0[28]) );
  INVX1 U9230 ( .A(n8315), .Y(N59) );
  AND2X1 U9231 ( .A(N58), .B(read_en[0]), .Y(rdata_0[29]) );
  INVX1 U9232 ( .A(n8316), .Y(N58) );
  AND2X1 U9233 ( .A(N57), .B(read_en[0]), .Y(rdata_0[30]) );
  INVX1 U9234 ( .A(n8317), .Y(N57) );
  AND2X1 U9235 ( .A(N56), .B(read_en[0]), .Y(rdata_0[31]) );
  INVX1 U9236 ( .A(n8318), .Y(N56) );
  AND2X1 U9237 ( .A(N55), .B(read_en[0]), .Y(rdata_0[32]) );
  INVX1 U9238 ( .A(n8319), .Y(N55) );
  AND2X1 U9239 ( .A(N54), .B(read_en[0]), .Y(rdata_0[33]) );
  INVX1 U9240 ( .A(n8320), .Y(N54) );
  AND2X1 U9241 ( .A(N53), .B(read_en[0]), .Y(rdata_0[34]) );
  INVX1 U9242 ( .A(n8321), .Y(N53) );
  AND2X1 U9243 ( .A(N52), .B(read_en[0]), .Y(rdata_0[35]) );
  INVX1 U9244 ( .A(n8322), .Y(N52) );
  AND2X1 U9245 ( .A(N51), .B(read_en[0]), .Y(rdata_0[36]) );
  INVX1 U9246 ( .A(n8323), .Y(N51) );
  AND2X1 U9247 ( .A(N50), .B(read_en[0]), .Y(rdata_0[37]) );
  INVX1 U9248 ( .A(n8324), .Y(N50) );
  AND2X1 U9249 ( .A(N49), .B(read_en[0]), .Y(rdata_0[38]) );
  INVX1 U9250 ( .A(n8325), .Y(N49) );
  AND2X1 U9251 ( .A(N48), .B(read_en[0]), .Y(rdata_0[39]) );
  INVX1 U9252 ( .A(n8326), .Y(N48) );
  AND2X1 U9253 ( .A(N47), .B(read_en[0]), .Y(rdata_0[40]) );
  INVX1 U9254 ( .A(n8327), .Y(N47) );
  AND2X1 U9255 ( .A(N46), .B(read_en[0]), .Y(rdata_0[41]) );
  INVX1 U9256 ( .A(n8328), .Y(N46) );
  AND2X1 U9257 ( .A(N45), .B(read_en[0]), .Y(rdata_0[42]) );
  INVX1 U9258 ( .A(n8329), .Y(N45) );
  AND2X1 U9259 ( .A(N44), .B(read_en[0]), .Y(rdata_0[43]) );
  INVX1 U9260 ( .A(n8330), .Y(N44) );
  AND2X1 U9261 ( .A(N43), .B(read_en[0]), .Y(rdata_0[44]) );
  INVX1 U9262 ( .A(n8331), .Y(N43) );
  AND2X1 U9263 ( .A(N42), .B(read_en[0]), .Y(rdata_0[45]) );
  INVX1 U9264 ( .A(n8332), .Y(N42) );
  AND2X1 U9265 ( .A(N41), .B(read_en[0]), .Y(rdata_0[46]) );
  INVX1 U9266 ( .A(n8333), .Y(N41) );
  AND2X1 U9267 ( .A(N40), .B(read_en[0]), .Y(rdata_0[47]) );
  INVX1 U9268 ( .A(n8334), .Y(N40) );
  AND2X1 U9269 ( .A(N39), .B(read_en[0]), .Y(rdata_0[48]) );
  INVX1 U9270 ( .A(n8335), .Y(N39) );
  AND2X1 U9271 ( .A(N38), .B(read_en[0]), .Y(rdata_0[49]) );
  INVX1 U9272 ( .A(n8336), .Y(N38) );
  AND2X1 U9273 ( .A(N37), .B(read_en[0]), .Y(rdata_0[50]) );
  INVX1 U9274 ( .A(n8337), .Y(N37) );
  AND2X1 U9275 ( .A(N36), .B(read_en[0]), .Y(rdata_0[51]) );
  INVX1 U9276 ( .A(n8338), .Y(N36) );
  AND2X1 U9277 ( .A(N35), .B(read_en[0]), .Y(rdata_0[52]) );
  INVX1 U9278 ( .A(n8339), .Y(N35) );
  AND2X1 U9279 ( .A(N34), .B(read_en[0]), .Y(rdata_0[53]) );
  INVX1 U9280 ( .A(n8340), .Y(N34) );
  AND2X1 U9281 ( .A(N33), .B(read_en[0]), .Y(rdata_0[54]) );
  INVX1 U9282 ( .A(n8341), .Y(N33) );
  AND2X1 U9283 ( .A(N32), .B(read_en[0]), .Y(rdata_0[55]) );
  INVX1 U9284 ( .A(n8342), .Y(N32) );
  AND2X1 U9285 ( .A(N31), .B(read_en[0]), .Y(rdata_0[56]) );
  INVX1 U9286 ( .A(n8343), .Y(N31) );
  AND2X1 U9287 ( .A(N30), .B(read_en[0]), .Y(rdata_0[57]) );
  INVX1 U9288 ( .A(n8344), .Y(N30) );
  AND2X1 U9289 ( .A(N29), .B(read_en[0]), .Y(rdata_0[58]) );
  INVX1 U9290 ( .A(n8345), .Y(N29) );
  AND2X1 U9291 ( .A(N28), .B(read_en[0]), .Y(rdata_0[59]) );
  INVX1 U9292 ( .A(n8346), .Y(N28) );
  AND2X1 U9293 ( .A(N27), .B(read_en[0]), .Y(rdata_0[60]) );
  INVX1 U9294 ( .A(n8347), .Y(N27) );
  AND2X1 U9295 ( .A(N26), .B(read_en[0]), .Y(rdata_0[61]) );
  INVX1 U9296 ( .A(n8348), .Y(N26) );
  AND2X1 U9297 ( .A(N25), .B(read_en[0]), .Y(rdata_0[62]) );
  INVX1 U9298 ( .A(n8349), .Y(N25) );
  AND2X1 U9299 ( .A(N24), .B(read_en[0]), .Y(rdata_0[63]) );
  INVX1 U9300 ( .A(n8350), .Y(N24) );
  INVX1 U9301 ( .A(waddr[4]), .Y(n10831) );
  INVX1 U9302 ( .A(waddr[3]), .Y(n10832) );
  MUX2X1 U9303 ( .B(n6368), .A(n6369), .S(n8472), .Y(n6367) );
  MUX2X1 U9304 ( .B(n6371), .A(n6372), .S(n8472), .Y(n6370) );
  MUX2X1 U9305 ( .B(n6374), .A(n6375), .S(n8472), .Y(n6373) );
  MUX2X1 U9306 ( .B(n6377), .A(n6378), .S(n8472), .Y(n6376) );
  MUX2X1 U9307 ( .B(n6380), .A(n6381), .S(N16), .Y(n6379) );
  MUX2X1 U9308 ( .B(n6383), .A(n6384), .S(n8472), .Y(n6382) );
  MUX2X1 U9309 ( .B(n6386), .A(n6387), .S(n8472), .Y(n6385) );
  MUX2X1 U9310 ( .B(n6389), .A(n6390), .S(n8472), .Y(n6388) );
  MUX2X1 U9311 ( .B(n6392), .A(n6393), .S(n8472), .Y(n6391) );
  MUX2X1 U9312 ( .B(n6395), .A(n6396), .S(N16), .Y(n6394) );
  MUX2X1 U9313 ( .B(n6398), .A(n6399), .S(n8473), .Y(n6397) );
  MUX2X1 U9314 ( .B(n6401), .A(n6402), .S(n8473), .Y(n6400) );
  MUX2X1 U9315 ( .B(n6404), .A(n6405), .S(n8473), .Y(n6403) );
  MUX2X1 U9316 ( .B(n6407), .A(n6408), .S(n8473), .Y(n6406) );
  MUX2X1 U9317 ( .B(n6410), .A(n6411), .S(N16), .Y(n6409) );
  MUX2X1 U9318 ( .B(n6413), .A(n6414), .S(n8473), .Y(n6412) );
  MUX2X1 U9319 ( .B(n6416), .A(n6417), .S(n8473), .Y(n6415) );
  MUX2X1 U9320 ( .B(n6419), .A(n6420), .S(n8473), .Y(n6418) );
  MUX2X1 U9321 ( .B(n6422), .A(n6423), .S(n8473), .Y(n6421) );
  MUX2X1 U9322 ( .B(n6425), .A(n6426), .S(N16), .Y(n6424) );
  MUX2X1 U9323 ( .B(n6428), .A(n6429), .S(n8473), .Y(n6427) );
  MUX2X1 U9324 ( .B(n6431), .A(n6432), .S(n8473), .Y(n6430) );
  MUX2X1 U9325 ( .B(n6434), .A(n6435), .S(n8473), .Y(n6433) );
  MUX2X1 U9326 ( .B(n6437), .A(n6438), .S(n8473), .Y(n6436) );
  MUX2X1 U9327 ( .B(n6440), .A(n6441), .S(N16), .Y(n6439) );
  MUX2X1 U9328 ( .B(n6443), .A(n6444), .S(n8474), .Y(n6442) );
  MUX2X1 U9329 ( .B(n6446), .A(n6447), .S(n8474), .Y(n6445) );
  MUX2X1 U9330 ( .B(n6449), .A(n6450), .S(n8474), .Y(n6448) );
  MUX2X1 U9331 ( .B(n6452), .A(n6453), .S(n8474), .Y(n6451) );
  MUX2X1 U9332 ( .B(n6455), .A(n6456), .S(N16), .Y(n6454) );
  MUX2X1 U9333 ( .B(n6458), .A(n6459), .S(n8474), .Y(n6457) );
  MUX2X1 U9334 ( .B(n6461), .A(n6462), .S(n8474), .Y(n6460) );
  MUX2X1 U9335 ( .B(n6464), .A(n6465), .S(n8474), .Y(n6463) );
  MUX2X1 U9336 ( .B(n6467), .A(n6468), .S(n8474), .Y(n6466) );
  MUX2X1 U9337 ( .B(n6470), .A(n6471), .S(N16), .Y(n6469) );
  MUX2X1 U9338 ( .B(n6473), .A(n6474), .S(n8474), .Y(n6472) );
  MUX2X1 U9339 ( .B(n6476), .A(n6477), .S(n8474), .Y(n6475) );
  MUX2X1 U9340 ( .B(n6479), .A(n6480), .S(n8474), .Y(n6478) );
  MUX2X1 U9341 ( .B(n6482), .A(n6483), .S(n8474), .Y(n6481) );
  MUX2X1 U9342 ( .B(n6485), .A(n6486), .S(N16), .Y(n6484) );
  MUX2X1 U9343 ( .B(n6488), .A(n6489), .S(n8475), .Y(n6487) );
  MUX2X1 U9344 ( .B(n6491), .A(n6492), .S(n8475), .Y(n6490) );
  MUX2X1 U9345 ( .B(n6494), .A(n6495), .S(n8475), .Y(n6493) );
  MUX2X1 U9346 ( .B(n6497), .A(n6498), .S(n8475), .Y(n6496) );
  MUX2X1 U9347 ( .B(n6500), .A(n6501), .S(N16), .Y(n6499) );
  MUX2X1 U9348 ( .B(n6503), .A(n6504), .S(n8475), .Y(n6502) );
  MUX2X1 U9349 ( .B(n6506), .A(n6507), .S(n8475), .Y(n6505) );
  MUX2X1 U9350 ( .B(n6509), .A(n6510), .S(n8475), .Y(n6508) );
  MUX2X1 U9351 ( .B(n6512), .A(n6513), .S(n8475), .Y(n6511) );
  MUX2X1 U9352 ( .B(n6515), .A(n6516), .S(N16), .Y(n6514) );
  MUX2X1 U9353 ( .B(n6518), .A(n6519), .S(n8475), .Y(n6517) );
  MUX2X1 U9354 ( .B(n6521), .A(n6522), .S(n8475), .Y(n6520) );
  MUX2X1 U9355 ( .B(n6524), .A(n6525), .S(n8475), .Y(n6523) );
  MUX2X1 U9356 ( .B(n6527), .A(n6528), .S(n8475), .Y(n6526) );
  MUX2X1 U9357 ( .B(n6530), .A(n6531), .S(N16), .Y(n6529) );
  MUX2X1 U9358 ( .B(n6533), .A(n6534), .S(n8476), .Y(n6532) );
  MUX2X1 U9359 ( .B(n6536), .A(n6537), .S(n8476), .Y(n6535) );
  MUX2X1 U9360 ( .B(n6539), .A(n6540), .S(n8476), .Y(n6538) );
  MUX2X1 U9361 ( .B(n6542), .A(n6543), .S(n8476), .Y(n6541) );
  MUX2X1 U9362 ( .B(n6545), .A(n6546), .S(N16), .Y(n6544) );
  MUX2X1 U9363 ( .B(n6548), .A(n6549), .S(n8476), .Y(n6547) );
  MUX2X1 U9364 ( .B(n6551), .A(n6552), .S(n8476), .Y(n6550) );
  MUX2X1 U9365 ( .B(n6554), .A(n6555), .S(n8476), .Y(n6553) );
  MUX2X1 U9366 ( .B(n6557), .A(n6558), .S(n8476), .Y(n6556) );
  MUX2X1 U9367 ( .B(n6560), .A(n6561), .S(N16), .Y(n6559) );
  MUX2X1 U9368 ( .B(n6563), .A(n6564), .S(n8476), .Y(n6562) );
  MUX2X1 U9369 ( .B(n6566), .A(n6567), .S(n8476), .Y(n6565) );
  MUX2X1 U9370 ( .B(n6569), .A(n6570), .S(n8476), .Y(n6568) );
  MUX2X1 U9371 ( .B(n6572), .A(n6573), .S(n8476), .Y(n6571) );
  MUX2X1 U9372 ( .B(n6575), .A(n6576), .S(N16), .Y(n6574) );
  MUX2X1 U9373 ( .B(n6578), .A(n6579), .S(n8477), .Y(n6577) );
  MUX2X1 U9374 ( .B(n6581), .A(n6582), .S(n8477), .Y(n6580) );
  MUX2X1 U9375 ( .B(n6584), .A(n6585), .S(n8477), .Y(n6583) );
  MUX2X1 U9376 ( .B(n6587), .A(n6588), .S(n8477), .Y(n6586) );
  MUX2X1 U9377 ( .B(n6590), .A(n6591), .S(N16), .Y(n6589) );
  MUX2X1 U9378 ( .B(n6593), .A(n6594), .S(n8477), .Y(n6592) );
  MUX2X1 U9379 ( .B(n6596), .A(n6597), .S(n8477), .Y(n6595) );
  MUX2X1 U9380 ( .B(n6599), .A(n6600), .S(n8477), .Y(n6598) );
  MUX2X1 U9381 ( .B(n6602), .A(n6603), .S(n8477), .Y(n6601) );
  MUX2X1 U9382 ( .B(n6605), .A(n6606), .S(N16), .Y(n6604) );
  MUX2X1 U9383 ( .B(n6608), .A(n6609), .S(n8477), .Y(n6607) );
  MUX2X1 U9384 ( .B(n6611), .A(n6612), .S(n8477), .Y(n6610) );
  MUX2X1 U9385 ( .B(n6614), .A(n6615), .S(n8477), .Y(n6613) );
  MUX2X1 U9386 ( .B(n6617), .A(n6618), .S(n8477), .Y(n6616) );
  MUX2X1 U9387 ( .B(n6620), .A(n6621), .S(N16), .Y(n6619) );
  MUX2X1 U9388 ( .B(n6623), .A(n6624), .S(n8478), .Y(n6622) );
  MUX2X1 U9389 ( .B(n6626), .A(n6627), .S(n8478), .Y(n6625) );
  MUX2X1 U9390 ( .B(n6629), .A(n6630), .S(n8478), .Y(n6628) );
  MUX2X1 U9391 ( .B(n6632), .A(n6633), .S(n8478), .Y(n6631) );
  MUX2X1 U9392 ( .B(n6635), .A(n6636), .S(N16), .Y(n6634) );
  MUX2X1 U9393 ( .B(n6638), .A(n6639), .S(n8478), .Y(n6637) );
  MUX2X1 U9394 ( .B(n6641), .A(n6642), .S(n8478), .Y(n6640) );
  MUX2X1 U9395 ( .B(n6644), .A(n6645), .S(n8478), .Y(n6643) );
  MUX2X1 U9396 ( .B(n6647), .A(n6648), .S(n8478), .Y(n6646) );
  MUX2X1 U9397 ( .B(n6650), .A(n6651), .S(N16), .Y(n6649) );
  MUX2X1 U9398 ( .B(n6653), .A(n6654), .S(n8478), .Y(n6652) );
  MUX2X1 U9399 ( .B(n6656), .A(n6657), .S(n8478), .Y(n6655) );
  MUX2X1 U9400 ( .B(n6659), .A(n6660), .S(n8478), .Y(n6658) );
  MUX2X1 U9401 ( .B(n6662), .A(n6663), .S(n8478), .Y(n6661) );
  MUX2X1 U9402 ( .B(n6665), .A(n6666), .S(N16), .Y(n6664) );
  MUX2X1 U9403 ( .B(n6668), .A(n6669), .S(n8479), .Y(n6667) );
  MUX2X1 U9404 ( .B(n6671), .A(n6672), .S(n8479), .Y(n6670) );
  MUX2X1 U9405 ( .B(n6674), .A(n6675), .S(n8479), .Y(n6673) );
  MUX2X1 U9406 ( .B(n6677), .A(n6678), .S(n8479), .Y(n6676) );
  MUX2X1 U9407 ( .B(n6680), .A(n6681), .S(N16), .Y(n6679) );
  MUX2X1 U9408 ( .B(n6683), .A(n6684), .S(n8479), .Y(n6682) );
  MUX2X1 U9409 ( .B(n6686), .A(n6687), .S(n8479), .Y(n6685) );
  MUX2X1 U9410 ( .B(n6689), .A(n6690), .S(n8479), .Y(n6688) );
  MUX2X1 U9411 ( .B(n6692), .A(n6693), .S(n8479), .Y(n6691) );
  MUX2X1 U9412 ( .B(n6695), .A(n6696), .S(N16), .Y(n6694) );
  MUX2X1 U9413 ( .B(n6698), .A(n6699), .S(n8479), .Y(n6697) );
  MUX2X1 U9414 ( .B(n6701), .A(n6702), .S(n8479), .Y(n6700) );
  MUX2X1 U9415 ( .B(n6704), .A(n6705), .S(n8479), .Y(n6703) );
  MUX2X1 U9416 ( .B(n6707), .A(n6708), .S(n8479), .Y(n6706) );
  MUX2X1 U9417 ( .B(n6710), .A(n6711), .S(N16), .Y(n6709) );
  MUX2X1 U9418 ( .B(n6713), .A(n6714), .S(n8480), .Y(n6712) );
  MUX2X1 U9419 ( .B(n6716), .A(n6717), .S(n8480), .Y(n6715) );
  MUX2X1 U9420 ( .B(n6719), .A(n6720), .S(n8480), .Y(n6718) );
  MUX2X1 U9421 ( .B(n6722), .A(n6723), .S(n8480), .Y(n6721) );
  MUX2X1 U9422 ( .B(n6725), .A(n6726), .S(N16), .Y(n6724) );
  MUX2X1 U9423 ( .B(n6728), .A(n6729), .S(n8480), .Y(n6727) );
  MUX2X1 U9424 ( .B(n6731), .A(n6732), .S(n8480), .Y(n6730) );
  MUX2X1 U9425 ( .B(n6734), .A(n6735), .S(n8480), .Y(n6733) );
  MUX2X1 U9426 ( .B(n6737), .A(n6738), .S(n8480), .Y(n6736) );
  MUX2X1 U9427 ( .B(n6740), .A(n6741), .S(N16), .Y(n6739) );
  MUX2X1 U9428 ( .B(n6743), .A(n6744), .S(n8480), .Y(n6742) );
  MUX2X1 U9429 ( .B(n6746), .A(n6747), .S(n8480), .Y(n6745) );
  MUX2X1 U9430 ( .B(n6749), .A(n6750), .S(n8480), .Y(n6748) );
  MUX2X1 U9431 ( .B(n6752), .A(n6753), .S(n8480), .Y(n6751) );
  MUX2X1 U9432 ( .B(n6755), .A(n6756), .S(N16), .Y(n6754) );
  MUX2X1 U9433 ( .B(n6758), .A(n6759), .S(n8481), .Y(n6757) );
  MUX2X1 U9434 ( .B(n6761), .A(n6762), .S(n8481), .Y(n6760) );
  MUX2X1 U9435 ( .B(n6764), .A(n6765), .S(n8481), .Y(n6763) );
  MUX2X1 U9436 ( .B(n6767), .A(n6768), .S(n8481), .Y(n6766) );
  MUX2X1 U9437 ( .B(n6770), .A(n6771), .S(N16), .Y(n6769) );
  MUX2X1 U9438 ( .B(n6773), .A(n6774), .S(n8481), .Y(n6772) );
  MUX2X1 U9439 ( .B(n6776), .A(n6777), .S(n8481), .Y(n6775) );
  MUX2X1 U9440 ( .B(n6779), .A(n6780), .S(n8481), .Y(n6778) );
  MUX2X1 U9441 ( .B(n6782), .A(n6783), .S(n8481), .Y(n6781) );
  MUX2X1 U9442 ( .B(n6785), .A(n6786), .S(N16), .Y(n6784) );
  MUX2X1 U9443 ( .B(n6788), .A(n6789), .S(n8481), .Y(n6787) );
  MUX2X1 U9444 ( .B(n6791), .A(n6792), .S(n8481), .Y(n6790) );
  MUX2X1 U9445 ( .B(n6794), .A(n6795), .S(n8481), .Y(n6793) );
  MUX2X1 U9446 ( .B(n6797), .A(n6798), .S(n8481), .Y(n6796) );
  MUX2X1 U9447 ( .B(n6800), .A(n6801), .S(N16), .Y(n6799) );
  MUX2X1 U9448 ( .B(n6803), .A(n6804), .S(n8482), .Y(n6802) );
  MUX2X1 U9449 ( .B(n6806), .A(n6807), .S(n8482), .Y(n6805) );
  MUX2X1 U9450 ( .B(n6809), .A(n6810), .S(n8482), .Y(n6808) );
  MUX2X1 U9451 ( .B(n6812), .A(n6813), .S(n8482), .Y(n6811) );
  MUX2X1 U9452 ( .B(n6815), .A(n6816), .S(N16), .Y(n6814) );
  MUX2X1 U9453 ( .B(n6818), .A(n6819), .S(n8482), .Y(n6817) );
  MUX2X1 U9454 ( .B(n6821), .A(n6822), .S(n8482), .Y(n6820) );
  MUX2X1 U9455 ( .B(n6824), .A(n6825), .S(n8482), .Y(n6823) );
  MUX2X1 U9456 ( .B(n6827), .A(n6828), .S(n8482), .Y(n6826) );
  MUX2X1 U9457 ( .B(n6830), .A(n6831), .S(N16), .Y(n6829) );
  MUX2X1 U9458 ( .B(n6833), .A(n6834), .S(n8482), .Y(n6832) );
  MUX2X1 U9459 ( .B(n6836), .A(n6837), .S(n8482), .Y(n6835) );
  MUX2X1 U9460 ( .B(n6839), .A(n6840), .S(n8482), .Y(n6838) );
  MUX2X1 U9461 ( .B(n6842), .A(n6843), .S(n8482), .Y(n6841) );
  MUX2X1 U9462 ( .B(n6845), .A(n6846), .S(N16), .Y(n6844) );
  MUX2X1 U9463 ( .B(n6848), .A(n6849), .S(n8483), .Y(n6847) );
  MUX2X1 U9464 ( .B(n6851), .A(n6852), .S(n8483), .Y(n6850) );
  MUX2X1 U9465 ( .B(n6854), .A(n6855), .S(n8483), .Y(n6853) );
  MUX2X1 U9466 ( .B(n6857), .A(n6858), .S(n8483), .Y(n6856) );
  MUX2X1 U9467 ( .B(n6860), .A(n6861), .S(N16), .Y(n6859) );
  MUX2X1 U9468 ( .B(n6863), .A(n6864), .S(n8483), .Y(n6862) );
  MUX2X1 U9469 ( .B(n6866), .A(n6867), .S(n8483), .Y(n6865) );
  MUX2X1 U9470 ( .B(n6869), .A(n6870), .S(n8483), .Y(n6868) );
  MUX2X1 U9471 ( .B(n6872), .A(n6873), .S(n8483), .Y(n6871) );
  MUX2X1 U9472 ( .B(n6875), .A(n6876), .S(N16), .Y(n6874) );
  MUX2X1 U9473 ( .B(n6878), .A(n6879), .S(n8483), .Y(n6877) );
  MUX2X1 U9474 ( .B(n6881), .A(n6882), .S(n8483), .Y(n6880) );
  MUX2X1 U9475 ( .B(n6884), .A(n6885), .S(n8483), .Y(n6883) );
  MUX2X1 U9476 ( .B(n6887), .A(n6888), .S(n8483), .Y(n6886) );
  MUX2X1 U9477 ( .B(n6890), .A(n6891), .S(N16), .Y(n6889) );
  MUX2X1 U9478 ( .B(n6893), .A(n6894), .S(n8484), .Y(n6892) );
  MUX2X1 U9479 ( .B(n6896), .A(n6897), .S(n8484), .Y(n6895) );
  MUX2X1 U9480 ( .B(n6899), .A(n6900), .S(n8484), .Y(n6898) );
  MUX2X1 U9481 ( .B(n6902), .A(n6903), .S(n8484), .Y(n6901) );
  MUX2X1 U9482 ( .B(n6905), .A(n6906), .S(N16), .Y(n6904) );
  MUX2X1 U9483 ( .B(n6908), .A(n6909), .S(n8484), .Y(n6907) );
  MUX2X1 U9484 ( .B(n6911), .A(n6912), .S(n8484), .Y(n6910) );
  MUX2X1 U9485 ( .B(n6914), .A(n6915), .S(n8484), .Y(n6913) );
  MUX2X1 U9486 ( .B(n6917), .A(n6918), .S(n8484), .Y(n6916) );
  MUX2X1 U9487 ( .B(n6920), .A(n6921), .S(N16), .Y(n6919) );
  MUX2X1 U9488 ( .B(n6923), .A(n6924), .S(n8484), .Y(n6922) );
  MUX2X1 U9489 ( .B(n6926), .A(n6927), .S(n8484), .Y(n6925) );
  MUX2X1 U9490 ( .B(n6929), .A(n6930), .S(n8484), .Y(n6928) );
  MUX2X1 U9491 ( .B(n6932), .A(n6933), .S(n8484), .Y(n6931) );
  MUX2X1 U9492 ( .B(n6935), .A(n6936), .S(N16), .Y(n6934) );
  MUX2X1 U9493 ( .B(n6938), .A(n6939), .S(n8485), .Y(n6937) );
  MUX2X1 U9494 ( .B(n6941), .A(n6942), .S(n8485), .Y(n6940) );
  MUX2X1 U9495 ( .B(n6944), .A(n6945), .S(n8485), .Y(n6943) );
  MUX2X1 U9496 ( .B(n6947), .A(n6948), .S(n8485), .Y(n6946) );
  MUX2X1 U9497 ( .B(n6950), .A(n6951), .S(N16), .Y(n6949) );
  MUX2X1 U9498 ( .B(n6953), .A(n6954), .S(n8485), .Y(n6952) );
  MUX2X1 U9499 ( .B(n6956), .A(n6957), .S(n8485), .Y(n6955) );
  MUX2X1 U9500 ( .B(n6959), .A(n6960), .S(n8485), .Y(n6958) );
  MUX2X1 U9501 ( .B(n6962), .A(n6963), .S(n8485), .Y(n6961) );
  MUX2X1 U9502 ( .B(n6965), .A(n6966), .S(N16), .Y(n6964) );
  MUX2X1 U9503 ( .B(n6968), .A(n6969), .S(n8485), .Y(n6967) );
  MUX2X1 U9504 ( .B(n6971), .A(n6972), .S(n8485), .Y(n6970) );
  MUX2X1 U9505 ( .B(n6974), .A(n6975), .S(n8485), .Y(n6973) );
  MUX2X1 U9506 ( .B(n6977), .A(n6978), .S(n8485), .Y(n6976) );
  MUX2X1 U9507 ( .B(n6980), .A(n6981), .S(N16), .Y(n6979) );
  MUX2X1 U9508 ( .B(n6983), .A(n6984), .S(n8486), .Y(n6982) );
  MUX2X1 U9509 ( .B(n6986), .A(n6987), .S(n8486), .Y(n6985) );
  MUX2X1 U9510 ( .B(n6989), .A(n6990), .S(n8486), .Y(n6988) );
  MUX2X1 U9511 ( .B(n6992), .A(n6993), .S(n8486), .Y(n6991) );
  MUX2X1 U9512 ( .B(n6995), .A(n6996), .S(N16), .Y(n6994) );
  MUX2X1 U9513 ( .B(n6998), .A(n6999), .S(n8486), .Y(n6997) );
  MUX2X1 U9514 ( .B(n7001), .A(n7002), .S(n8486), .Y(n7000) );
  MUX2X1 U9515 ( .B(n7004), .A(n7005), .S(n8486), .Y(n7003) );
  MUX2X1 U9516 ( .B(n7007), .A(n7008), .S(n8486), .Y(n7006) );
  MUX2X1 U9517 ( .B(n7010), .A(n7011), .S(N16), .Y(n7009) );
  MUX2X1 U9518 ( .B(n7013), .A(n7014), .S(n8486), .Y(n7012) );
  MUX2X1 U9519 ( .B(n7016), .A(n7017), .S(n8486), .Y(n7015) );
  MUX2X1 U9520 ( .B(n7019), .A(n7020), .S(n8486), .Y(n7018) );
  MUX2X1 U9521 ( .B(n7022), .A(n7023), .S(n8486), .Y(n7021) );
  MUX2X1 U9522 ( .B(n7025), .A(n7026), .S(N16), .Y(n7024) );
  MUX2X1 U9523 ( .B(n7028), .A(n7029), .S(n8487), .Y(n7027) );
  MUX2X1 U9524 ( .B(n7031), .A(n7032), .S(n8487), .Y(n7030) );
  MUX2X1 U9525 ( .B(n7034), .A(n7035), .S(n8487), .Y(n7033) );
  MUX2X1 U9526 ( .B(n7037), .A(n7038), .S(n8487), .Y(n7036) );
  MUX2X1 U9527 ( .B(n7040), .A(n7041), .S(N16), .Y(n7039) );
  MUX2X1 U9528 ( .B(n7043), .A(n7044), .S(n8487), .Y(n7042) );
  MUX2X1 U9529 ( .B(n7046), .A(n7047), .S(n8487), .Y(n7045) );
  MUX2X1 U9530 ( .B(n7049), .A(n7050), .S(n8487), .Y(n7048) );
  MUX2X1 U9531 ( .B(n7052), .A(n7053), .S(n8487), .Y(n7051) );
  MUX2X1 U9532 ( .B(n7055), .A(n7056), .S(N16), .Y(n7054) );
  MUX2X1 U9533 ( .B(n7058), .A(n7059), .S(n8487), .Y(n7057) );
  MUX2X1 U9534 ( .B(n7061), .A(n7062), .S(n8487), .Y(n7060) );
  MUX2X1 U9535 ( .B(n7064), .A(n7065), .S(n8487), .Y(n7063) );
  MUX2X1 U9536 ( .B(n7067), .A(n7068), .S(n8487), .Y(n7066) );
  MUX2X1 U9537 ( .B(n7070), .A(n7071), .S(N16), .Y(n7069) );
  MUX2X1 U9538 ( .B(n7073), .A(n7074), .S(n8488), .Y(n7072) );
  MUX2X1 U9539 ( .B(n7076), .A(n7077), .S(n8488), .Y(n7075) );
  MUX2X1 U9540 ( .B(n7079), .A(n7080), .S(n8488), .Y(n7078) );
  MUX2X1 U9541 ( .B(n7082), .A(n7083), .S(n8488), .Y(n7081) );
  MUX2X1 U9542 ( .B(n7085), .A(n7086), .S(N16), .Y(n7084) );
  MUX2X1 U9543 ( .B(n7088), .A(n7089), .S(n8488), .Y(n7087) );
  MUX2X1 U9544 ( .B(n7091), .A(n7092), .S(n8488), .Y(n7090) );
  MUX2X1 U9545 ( .B(n7094), .A(n7095), .S(n8488), .Y(n7093) );
  MUX2X1 U9546 ( .B(n7097), .A(n7098), .S(n8488), .Y(n7096) );
  MUX2X1 U9547 ( .B(n7100), .A(n7101), .S(N16), .Y(n7099) );
  MUX2X1 U9548 ( .B(n7103), .A(n7104), .S(n8488), .Y(n7102) );
  MUX2X1 U9549 ( .B(n7106), .A(n7107), .S(n8488), .Y(n7105) );
  MUX2X1 U9550 ( .B(n7109), .A(n7110), .S(n8488), .Y(n7108) );
  MUX2X1 U9551 ( .B(n7112), .A(n7113), .S(n8488), .Y(n7111) );
  MUX2X1 U9552 ( .B(n7115), .A(n7116), .S(N16), .Y(n7114) );
  MUX2X1 U9553 ( .B(n7118), .A(n7119), .S(n8489), .Y(n7117) );
  MUX2X1 U9554 ( .B(n7121), .A(n7122), .S(n8489), .Y(n7120) );
  MUX2X1 U9555 ( .B(n7124), .A(n7125), .S(n8489), .Y(n7123) );
  MUX2X1 U9556 ( .B(n7127), .A(n7128), .S(n8489), .Y(n7126) );
  MUX2X1 U9557 ( .B(n7130), .A(n7131), .S(N16), .Y(n7129) );
  MUX2X1 U9558 ( .B(n7133), .A(n7134), .S(n8489), .Y(n7132) );
  MUX2X1 U9559 ( .B(n7136), .A(n7137), .S(n8489), .Y(n7135) );
  MUX2X1 U9560 ( .B(n7139), .A(n7140), .S(n8489), .Y(n7138) );
  MUX2X1 U9561 ( .B(n7142), .A(n7143), .S(n8489), .Y(n7141) );
  MUX2X1 U9562 ( .B(n7145), .A(n7146), .S(N16), .Y(n7144) );
  MUX2X1 U9563 ( .B(n7148), .A(n7149), .S(n8489), .Y(n7147) );
  MUX2X1 U9564 ( .B(n7151), .A(n7152), .S(n8489), .Y(n7150) );
  MUX2X1 U9565 ( .B(n7154), .A(n7155), .S(n8489), .Y(n7153) );
  MUX2X1 U9566 ( .B(n7157), .A(n7158), .S(n8489), .Y(n7156) );
  MUX2X1 U9567 ( .B(n7160), .A(n7161), .S(N16), .Y(n7159) );
  MUX2X1 U9568 ( .B(n7163), .A(n7164), .S(n8490), .Y(n7162) );
  MUX2X1 U9569 ( .B(n7166), .A(n7167), .S(n8490), .Y(n7165) );
  MUX2X1 U9570 ( .B(n7169), .A(n7170), .S(n8490), .Y(n7168) );
  MUX2X1 U9571 ( .B(n7172), .A(n7173), .S(n8490), .Y(n7171) );
  MUX2X1 U9572 ( .B(n7175), .A(n7176), .S(N16), .Y(n7174) );
  MUX2X1 U9573 ( .B(n7178), .A(n7179), .S(n8490), .Y(n7177) );
  MUX2X1 U9574 ( .B(n7181), .A(n7182), .S(n8490), .Y(n7180) );
  MUX2X1 U9575 ( .B(n7184), .A(n7185), .S(n8490), .Y(n7183) );
  MUX2X1 U9576 ( .B(n7187), .A(n7188), .S(n8490), .Y(n7186) );
  MUX2X1 U9577 ( .B(n7190), .A(n7191), .S(N16), .Y(n7189) );
  MUX2X1 U9578 ( .B(n7193), .A(n7194), .S(n8490), .Y(n7192) );
  MUX2X1 U9579 ( .B(n7196), .A(n7197), .S(n8490), .Y(n7195) );
  MUX2X1 U9580 ( .B(n7199), .A(n7200), .S(n8490), .Y(n7198) );
  MUX2X1 U9581 ( .B(n7202), .A(n7203), .S(n8490), .Y(n7201) );
  MUX2X1 U9582 ( .B(n7205), .A(n7206), .S(N16), .Y(n7204) );
  MUX2X1 U9583 ( .B(n7208), .A(n7209), .S(n8491), .Y(n7207) );
  MUX2X1 U9584 ( .B(n7211), .A(n7212), .S(n8491), .Y(n7210) );
  MUX2X1 U9585 ( .B(n7214), .A(n7215), .S(n8491), .Y(n7213) );
  MUX2X1 U9586 ( .B(n7217), .A(n7218), .S(n8491), .Y(n7216) );
  MUX2X1 U9587 ( .B(n7220), .A(n7221), .S(N16), .Y(n7219) );
  MUX2X1 U9588 ( .B(n7223), .A(n7224), .S(n8491), .Y(n7222) );
  MUX2X1 U9589 ( .B(n7226), .A(n7227), .S(n8491), .Y(n7225) );
  MUX2X1 U9590 ( .B(n7229), .A(n7230), .S(n8491), .Y(n7228) );
  MUX2X1 U9591 ( .B(n7232), .A(n7233), .S(n8491), .Y(n7231) );
  MUX2X1 U9592 ( .B(n7235), .A(n7236), .S(N16), .Y(n7234) );
  MUX2X1 U9593 ( .B(n7238), .A(n7239), .S(n8491), .Y(n7237) );
  MUX2X1 U9594 ( .B(n7241), .A(n7242), .S(n8491), .Y(n7240) );
  MUX2X1 U9595 ( .B(n7244), .A(n7245), .S(n8491), .Y(n7243) );
  MUX2X1 U9596 ( .B(n7247), .A(n7248), .S(n8491), .Y(n7246) );
  MUX2X1 U9597 ( .B(n7250), .A(n7251), .S(N16), .Y(n7249) );
  MUX2X1 U9598 ( .B(n7253), .A(n7254), .S(n8492), .Y(n7252) );
  MUX2X1 U9599 ( .B(n7256), .A(n7257), .S(n8492), .Y(n7255) );
  MUX2X1 U9600 ( .B(n7259), .A(n7260), .S(n8492), .Y(n7258) );
  MUX2X1 U9601 ( .B(n7262), .A(n7263), .S(n8492), .Y(n7261) );
  MUX2X1 U9602 ( .B(n7265), .A(n7266), .S(N16), .Y(n7264) );
  MUX2X1 U9603 ( .B(n7268), .A(n7269), .S(n8492), .Y(n7267) );
  MUX2X1 U9604 ( .B(n7271), .A(n7272), .S(n8492), .Y(n7270) );
  MUX2X1 U9605 ( .B(n7274), .A(n7275), .S(n8492), .Y(n7273) );
  MUX2X1 U9606 ( .B(n7277), .A(n7278), .S(n8492), .Y(n7276) );
  MUX2X1 U9607 ( .B(n7280), .A(n7281), .S(N16), .Y(n7279) );
  MUX2X1 U9608 ( .B(n7283), .A(n7284), .S(n8492), .Y(n7282) );
  MUX2X1 U9609 ( .B(n7286), .A(n7287), .S(n8492), .Y(n7285) );
  MUX2X1 U9610 ( .B(n7289), .A(n7290), .S(n8492), .Y(n7288) );
  MUX2X1 U9611 ( .B(n7292), .A(n7293), .S(n8492), .Y(n7291) );
  MUX2X1 U9612 ( .B(n7295), .A(n7296), .S(N16), .Y(n7294) );
  MUX2X1 U9613 ( .B(n7298), .A(n7299), .S(n8493), .Y(n7297) );
  MUX2X1 U9614 ( .B(n7301), .A(n7302), .S(n8493), .Y(n7300) );
  MUX2X1 U9615 ( .B(n7304), .A(n7305), .S(n8493), .Y(n7303) );
  MUX2X1 U9616 ( .B(n7307), .A(n7308), .S(n8493), .Y(n7306) );
  MUX2X1 U9617 ( .B(n7310), .A(n7311), .S(N16), .Y(n7309) );
  MUX2X1 U9618 ( .B(n7313), .A(n7314), .S(n8493), .Y(n7312) );
  MUX2X1 U9619 ( .B(n7316), .A(n7317), .S(n8493), .Y(n7315) );
  MUX2X1 U9620 ( .B(n7319), .A(n7320), .S(n8493), .Y(n7318) );
  MUX2X1 U9621 ( .B(n7322), .A(n7323), .S(n8493), .Y(n7321) );
  MUX2X1 U9622 ( .B(n7325), .A(n7326), .S(N16), .Y(n7324) );
  MUX2X1 U9623 ( .B(n7328), .A(n7329), .S(n8493), .Y(n7327) );
  MUX2X1 U9624 ( .B(n7331), .A(n7332), .S(n8493), .Y(n7330) );
  MUX2X1 U9625 ( .B(n7334), .A(n7335), .S(n8493), .Y(n7333) );
  MUX2X1 U9626 ( .B(n7337), .A(n7338), .S(n8493), .Y(n7336) );
  MUX2X1 U9627 ( .B(n7340), .A(n7341), .S(N16), .Y(n7339) );
  MUX2X1 U9628 ( .B(n7343), .A(n7344), .S(n8494), .Y(n7342) );
  MUX2X1 U9629 ( .B(n7346), .A(n7347), .S(n8494), .Y(n7345) );
  MUX2X1 U9630 ( .B(n7349), .A(n7350), .S(n8494), .Y(n7348) );
  MUX2X1 U9631 ( .B(n7352), .A(n7353), .S(n8494), .Y(n7351) );
  MUX2X1 U9632 ( .B(n7355), .A(n7356), .S(N16), .Y(n7354) );
  MUX2X1 U9633 ( .B(n7358), .A(n7359), .S(n8494), .Y(n7357) );
  MUX2X1 U9634 ( .B(n7361), .A(n7362), .S(n8494), .Y(n7360) );
  MUX2X1 U9635 ( .B(n7364), .A(n7365), .S(n8494), .Y(n7363) );
  MUX2X1 U9636 ( .B(n7367), .A(n7368), .S(n8494), .Y(n7366) );
  MUX2X1 U9637 ( .B(n7370), .A(n7371), .S(N16), .Y(n7369) );
  MUX2X1 U9638 ( .B(n7373), .A(n7374), .S(n8494), .Y(n7372) );
  MUX2X1 U9639 ( .B(n7376), .A(n7377), .S(n8494), .Y(n7375) );
  MUX2X1 U9640 ( .B(n7379), .A(n7380), .S(n8494), .Y(n7378) );
  MUX2X1 U9641 ( .B(n7382), .A(n7383), .S(n8494), .Y(n7381) );
  MUX2X1 U9642 ( .B(n7385), .A(n7386), .S(N16), .Y(n7384) );
  MUX2X1 U9643 ( .B(n7388), .A(n7389), .S(n8495), .Y(n7387) );
  MUX2X1 U9644 ( .B(n7391), .A(n7392), .S(n8495), .Y(n7390) );
  MUX2X1 U9645 ( .B(n7394), .A(n7395), .S(n8495), .Y(n7393) );
  MUX2X1 U9646 ( .B(n7397), .A(n7398), .S(n8495), .Y(n7396) );
  MUX2X1 U9647 ( .B(n7400), .A(n7401), .S(N16), .Y(n7399) );
  MUX2X1 U9648 ( .B(n7403), .A(n7404), .S(n8495), .Y(n7402) );
  MUX2X1 U9649 ( .B(n7406), .A(n7407), .S(n8495), .Y(n7405) );
  MUX2X1 U9650 ( .B(n7409), .A(n7410), .S(n8495), .Y(n7408) );
  MUX2X1 U9651 ( .B(n7412), .A(n7413), .S(n8495), .Y(n7411) );
  MUX2X1 U9652 ( .B(n7415), .A(n7416), .S(N16), .Y(n7414) );
  MUX2X1 U9653 ( .B(n7418), .A(n7419), .S(n8495), .Y(n7417) );
  MUX2X1 U9654 ( .B(n7421), .A(n7422), .S(n8495), .Y(n7420) );
  MUX2X1 U9655 ( .B(n7424), .A(n7425), .S(n8495), .Y(n7423) );
  MUX2X1 U9656 ( .B(n7427), .A(n7428), .S(n8495), .Y(n7426) );
  MUX2X1 U9657 ( .B(n7430), .A(n7431), .S(N16), .Y(n7429) );
  MUX2X1 U9658 ( .B(n7433), .A(n7434), .S(n8496), .Y(n7432) );
  MUX2X1 U9659 ( .B(n7436), .A(n7437), .S(n8496), .Y(n7435) );
  MUX2X1 U9660 ( .B(n7439), .A(n7440), .S(n8496), .Y(n7438) );
  MUX2X1 U9661 ( .B(n7442), .A(n7443), .S(n8496), .Y(n7441) );
  MUX2X1 U9662 ( .B(n7445), .A(n7446), .S(N16), .Y(n7444) );
  MUX2X1 U9663 ( .B(n7448), .A(n7449), .S(n8496), .Y(n7447) );
  MUX2X1 U9664 ( .B(n7451), .A(n7452), .S(n8496), .Y(n7450) );
  MUX2X1 U9665 ( .B(n7454), .A(n7455), .S(n8496), .Y(n7453) );
  MUX2X1 U9666 ( .B(n7457), .A(n7458), .S(n8496), .Y(n7456) );
  MUX2X1 U9667 ( .B(n7460), .A(n7461), .S(N16), .Y(n7459) );
  MUX2X1 U9668 ( .B(n7463), .A(n7464), .S(n8496), .Y(n7462) );
  MUX2X1 U9669 ( .B(n7466), .A(n7467), .S(n8496), .Y(n7465) );
  MUX2X1 U9670 ( .B(n7469), .A(n7470), .S(n8496), .Y(n7468) );
  MUX2X1 U9671 ( .B(n7472), .A(n7473), .S(n8496), .Y(n7471) );
  MUX2X1 U9672 ( .B(n7475), .A(n7476), .S(N16), .Y(n7474) );
  MUX2X1 U9673 ( .B(n7478), .A(n7479), .S(n8497), .Y(n7477) );
  MUX2X1 U9674 ( .B(n7481), .A(n7482), .S(n8497), .Y(n7480) );
  MUX2X1 U9675 ( .B(n7484), .A(n7485), .S(n8497), .Y(n7483) );
  MUX2X1 U9676 ( .B(n7487), .A(n7488), .S(n8497), .Y(n7486) );
  MUX2X1 U9677 ( .B(n7490), .A(n7491), .S(N16), .Y(n7489) );
  MUX2X1 U9678 ( .B(n7493), .A(n7494), .S(n8497), .Y(n7492) );
  MUX2X1 U9679 ( .B(n7496), .A(n7497), .S(n8497), .Y(n7495) );
  MUX2X1 U9680 ( .B(n7499), .A(n7500), .S(n8497), .Y(n7498) );
  MUX2X1 U9681 ( .B(n7502), .A(n7503), .S(n8497), .Y(n7501) );
  MUX2X1 U9682 ( .B(n7505), .A(n7506), .S(N16), .Y(n7504) );
  MUX2X1 U9683 ( .B(n7508), .A(n7509), .S(n8497), .Y(n7507) );
  MUX2X1 U9684 ( .B(n7511), .A(n7512), .S(n8497), .Y(n7510) );
  MUX2X1 U9685 ( .B(n7514), .A(n7515), .S(n8497), .Y(n7513) );
  MUX2X1 U9686 ( .B(n7517), .A(n7518), .S(n8497), .Y(n7516) );
  MUX2X1 U9687 ( .B(n7520), .A(n7521), .S(N16), .Y(n7519) );
  MUX2X1 U9688 ( .B(n7523), .A(n7524), .S(n8498), .Y(n7522) );
  MUX2X1 U9689 ( .B(n7526), .A(n7527), .S(n8498), .Y(n7525) );
  MUX2X1 U9690 ( .B(n7529), .A(n7530), .S(n8498), .Y(n7528) );
  MUX2X1 U9691 ( .B(n7532), .A(n7533), .S(n8498), .Y(n7531) );
  MUX2X1 U9692 ( .B(n7535), .A(n7536), .S(N16), .Y(n7534) );
  MUX2X1 U9693 ( .B(n7538), .A(n7539), .S(n8498), .Y(n7537) );
  MUX2X1 U9694 ( .B(n7541), .A(n7542), .S(n8498), .Y(n7540) );
  MUX2X1 U9695 ( .B(n7544), .A(n7545), .S(n8498), .Y(n7543) );
  MUX2X1 U9696 ( .B(n7547), .A(n7548), .S(n8498), .Y(n7546) );
  MUX2X1 U9697 ( .B(n7550), .A(n7551), .S(N16), .Y(n7549) );
  MUX2X1 U9698 ( .B(n7553), .A(n7554), .S(n8498), .Y(n7552) );
  MUX2X1 U9699 ( .B(n7556), .A(n7557), .S(n8498), .Y(n7555) );
  MUX2X1 U9700 ( .B(n7559), .A(n7560), .S(n8498), .Y(n7558) );
  MUX2X1 U9701 ( .B(n7562), .A(n7563), .S(n8498), .Y(n7561) );
  MUX2X1 U9702 ( .B(n7565), .A(n7566), .S(N16), .Y(n7564) );
  MUX2X1 U9703 ( .B(n7568), .A(n7569), .S(n8499), .Y(n7567) );
  MUX2X1 U9704 ( .B(n7571), .A(n7572), .S(n8499), .Y(n7570) );
  MUX2X1 U9705 ( .B(n7574), .A(n7575), .S(n8499), .Y(n7573) );
  MUX2X1 U9706 ( .B(n7577), .A(n7578), .S(n8499), .Y(n7576) );
  MUX2X1 U9707 ( .B(n7580), .A(n7581), .S(N16), .Y(n7579) );
  MUX2X1 U9708 ( .B(n7583), .A(n7584), .S(n8499), .Y(n7582) );
  MUX2X1 U9709 ( .B(n7586), .A(n7587), .S(n8499), .Y(n7585) );
  MUX2X1 U9710 ( .B(n7589), .A(n7590), .S(n8499), .Y(n7588) );
  MUX2X1 U9711 ( .B(n7592), .A(n7593), .S(n8499), .Y(n7591) );
  MUX2X1 U9712 ( .B(n7595), .A(n7596), .S(N16), .Y(n7594) );
  MUX2X1 U9713 ( .B(n7598), .A(n7599), .S(n8499), .Y(n7597) );
  MUX2X1 U9714 ( .B(n7601), .A(n7602), .S(n8499), .Y(n7600) );
  MUX2X1 U9715 ( .B(n7604), .A(n7605), .S(n8499), .Y(n7603) );
  MUX2X1 U9716 ( .B(n7607), .A(n7608), .S(n8499), .Y(n7606) );
  MUX2X1 U9717 ( .B(n7610), .A(n7611), .S(N16), .Y(n7609) );
  MUX2X1 U9718 ( .B(n7613), .A(n7614), .S(n8500), .Y(n7612) );
  MUX2X1 U9719 ( .B(n7616), .A(n7617), .S(n8500), .Y(n7615) );
  MUX2X1 U9720 ( .B(n7619), .A(n7620), .S(n8500), .Y(n7618) );
  MUX2X1 U9721 ( .B(n7622), .A(n7623), .S(n8500), .Y(n7621) );
  MUX2X1 U9722 ( .B(n7625), .A(n7626), .S(N16), .Y(n7624) );
  MUX2X1 U9723 ( .B(n7628), .A(n7629), .S(n8500), .Y(n7627) );
  MUX2X1 U9724 ( .B(n7631), .A(n7632), .S(n8500), .Y(n7630) );
  MUX2X1 U9725 ( .B(n7634), .A(n7635), .S(n8500), .Y(n7633) );
  MUX2X1 U9726 ( .B(n7637), .A(n7638), .S(n8500), .Y(n7636) );
  MUX2X1 U9727 ( .B(n7640), .A(n7641), .S(N16), .Y(n7639) );
  MUX2X1 U9728 ( .B(n7643), .A(n7644), .S(n8500), .Y(n7642) );
  MUX2X1 U9729 ( .B(n7646), .A(n7647), .S(n8500), .Y(n7645) );
  MUX2X1 U9730 ( .B(n7649), .A(n7650), .S(n8500), .Y(n7648) );
  MUX2X1 U9731 ( .B(n7652), .A(n7653), .S(n8500), .Y(n7651) );
  MUX2X1 U9732 ( .B(n7655), .A(n7656), .S(N16), .Y(n7654) );
  MUX2X1 U9733 ( .B(n7658), .A(n7659), .S(n8501), .Y(n7657) );
  MUX2X1 U9734 ( .B(n7661), .A(n7662), .S(n8501), .Y(n7660) );
  MUX2X1 U9735 ( .B(n7664), .A(n7665), .S(n8501), .Y(n7663) );
  MUX2X1 U9736 ( .B(n7667), .A(n7668), .S(n8501), .Y(n7666) );
  MUX2X1 U9737 ( .B(n7670), .A(n7671), .S(N16), .Y(n7669) );
  MUX2X1 U9738 ( .B(n7673), .A(n7674), .S(n8501), .Y(n7672) );
  MUX2X1 U9739 ( .B(n7676), .A(n7677), .S(n8501), .Y(n7675) );
  MUX2X1 U9740 ( .B(n7679), .A(n7680), .S(n8501), .Y(n7678) );
  MUX2X1 U9741 ( .B(n7682), .A(n7683), .S(n8501), .Y(n7681) );
  MUX2X1 U9742 ( .B(n7685), .A(n7686), .S(N16), .Y(n7684) );
  MUX2X1 U9743 ( .B(n7688), .A(n7689), .S(n8501), .Y(n7687) );
  MUX2X1 U9744 ( .B(n7691), .A(n7692), .S(n8501), .Y(n7690) );
  MUX2X1 U9745 ( .B(n7694), .A(n7695), .S(n8501), .Y(n7693) );
  MUX2X1 U9746 ( .B(n7697), .A(n7698), .S(n8501), .Y(n7696) );
  MUX2X1 U9747 ( .B(n7700), .A(n7701), .S(N16), .Y(n7699) );
  MUX2X1 U9748 ( .B(n7703), .A(n7704), .S(n8502), .Y(n7702) );
  MUX2X1 U9749 ( .B(n7706), .A(n7707), .S(n8502), .Y(n7705) );
  MUX2X1 U9750 ( .B(n7709), .A(n7710), .S(n8502), .Y(n7708) );
  MUX2X1 U9751 ( .B(n7712), .A(n7713), .S(n8502), .Y(n7711) );
  MUX2X1 U9752 ( .B(n7715), .A(n7716), .S(N16), .Y(n7714) );
  MUX2X1 U9753 ( .B(n7718), .A(n7719), .S(n8502), .Y(n7717) );
  MUX2X1 U9754 ( .B(n7721), .A(n7722), .S(n8502), .Y(n7720) );
  MUX2X1 U9755 ( .B(n7724), .A(n7725), .S(n8502), .Y(n7723) );
  MUX2X1 U9756 ( .B(n7727), .A(n7728), .S(n8502), .Y(n7726) );
  MUX2X1 U9757 ( .B(n7730), .A(n7731), .S(N16), .Y(n7729) );
  MUX2X1 U9758 ( .B(n7733), .A(n7734), .S(n8502), .Y(n7732) );
  MUX2X1 U9759 ( .B(n7736), .A(n7737), .S(n8502), .Y(n7735) );
  MUX2X1 U9760 ( .B(n7739), .A(n7740), .S(n8502), .Y(n7738) );
  MUX2X1 U9761 ( .B(n7742), .A(n7743), .S(n8502), .Y(n7741) );
  MUX2X1 U9762 ( .B(n7745), .A(n7746), .S(N16), .Y(n7744) );
  MUX2X1 U9763 ( .B(n7748), .A(n7749), .S(n8503), .Y(n7747) );
  MUX2X1 U9764 ( .B(n7751), .A(n7752), .S(n8503), .Y(n7750) );
  MUX2X1 U9765 ( .B(n7754), .A(n7755), .S(n8503), .Y(n7753) );
  MUX2X1 U9766 ( .B(n7757), .A(n7758), .S(n8503), .Y(n7756) );
  MUX2X1 U9767 ( .B(n7760), .A(n7761), .S(N16), .Y(n7759) );
  MUX2X1 U9768 ( .B(n7763), .A(n7764), .S(n8503), .Y(n7762) );
  MUX2X1 U9769 ( .B(n7766), .A(n7767), .S(n8503), .Y(n7765) );
  MUX2X1 U9770 ( .B(n7769), .A(n7770), .S(n8503), .Y(n7768) );
  MUX2X1 U9771 ( .B(n7772), .A(n7773), .S(n8503), .Y(n7771) );
  MUX2X1 U9772 ( .B(n7775), .A(n7776), .S(N16), .Y(n7774) );
  MUX2X1 U9773 ( .B(n7778), .A(n7779), .S(n8503), .Y(n7777) );
  MUX2X1 U9774 ( .B(n7781), .A(n7782), .S(n8503), .Y(n7780) );
  MUX2X1 U9775 ( .B(n7784), .A(n7785), .S(n8503), .Y(n7783) );
  MUX2X1 U9776 ( .B(n7787), .A(n7788), .S(n8503), .Y(n7786) );
  MUX2X1 U9777 ( .B(n7790), .A(n7791), .S(N16), .Y(n7789) );
  MUX2X1 U9778 ( .B(n7793), .A(n7794), .S(n8504), .Y(n7792) );
  MUX2X1 U9779 ( .B(n7796), .A(n7797), .S(n8504), .Y(n7795) );
  MUX2X1 U9780 ( .B(n7799), .A(n7800), .S(n8504), .Y(n7798) );
  MUX2X1 U9781 ( .B(n7802), .A(n7803), .S(n8504), .Y(n7801) );
  MUX2X1 U9782 ( .B(n7805), .A(n7806), .S(N16), .Y(n7804) );
  MUX2X1 U9783 ( .B(n7808), .A(n7809), .S(n8504), .Y(n7807) );
  MUX2X1 U9784 ( .B(n7811), .A(n7812), .S(n8504), .Y(n7810) );
  MUX2X1 U9785 ( .B(n7814), .A(n7815), .S(n8504), .Y(n7813) );
  MUX2X1 U9786 ( .B(n7817), .A(n7818), .S(n8504), .Y(n7816) );
  MUX2X1 U9787 ( .B(n7820), .A(n7821), .S(N16), .Y(n7819) );
  MUX2X1 U9788 ( .B(n7823), .A(n7824), .S(n8504), .Y(n7822) );
  MUX2X1 U9789 ( .B(n7826), .A(n7827), .S(n8504), .Y(n7825) );
  MUX2X1 U9790 ( .B(n7829), .A(n7830), .S(n8504), .Y(n7828) );
  MUX2X1 U9791 ( .B(n7832), .A(n7833), .S(n8504), .Y(n7831) );
  MUX2X1 U9792 ( .B(n7835), .A(n7836), .S(N16), .Y(n7834) );
  MUX2X1 U9793 ( .B(n7838), .A(n7839), .S(n8505), .Y(n7837) );
  MUX2X1 U9794 ( .B(n7841), .A(n7842), .S(n8505), .Y(n7840) );
  MUX2X1 U9795 ( .B(n7844), .A(n7845), .S(n8505), .Y(n7843) );
  MUX2X1 U9796 ( .B(n7847), .A(n7848), .S(n8505), .Y(n7846) );
  MUX2X1 U9797 ( .B(n7850), .A(n7851), .S(N16), .Y(n7849) );
  MUX2X1 U9798 ( .B(n7853), .A(n7854), .S(n8505), .Y(n7852) );
  MUX2X1 U9799 ( .B(n7856), .A(n7857), .S(n8505), .Y(n7855) );
  MUX2X1 U9800 ( .B(n7859), .A(n7860), .S(n8505), .Y(n7858) );
  MUX2X1 U9801 ( .B(n7862), .A(n7863), .S(n8505), .Y(n7861) );
  MUX2X1 U9802 ( .B(n7865), .A(n7866), .S(N16), .Y(n7864) );
  MUX2X1 U9803 ( .B(n7868), .A(n7869), .S(n8505), .Y(n7867) );
  MUX2X1 U9804 ( .B(n7871), .A(n7872), .S(n8505), .Y(n7870) );
  MUX2X1 U9805 ( .B(n7874), .A(n7875), .S(n8505), .Y(n7873) );
  MUX2X1 U9806 ( .B(n7877), .A(n7878), .S(n8505), .Y(n7876) );
  MUX2X1 U9807 ( .B(n7880), .A(n7881), .S(N16), .Y(n7879) );
  MUX2X1 U9808 ( .B(n7883), .A(n7884), .S(n8506), .Y(n7882) );
  MUX2X1 U9809 ( .B(n7886), .A(n7887), .S(n8506), .Y(n7885) );
  MUX2X1 U9810 ( .B(n7889), .A(n7890), .S(n8506), .Y(n7888) );
  MUX2X1 U9811 ( .B(n7892), .A(n7893), .S(n8506), .Y(n7891) );
  MUX2X1 U9812 ( .B(n7895), .A(n7896), .S(N16), .Y(n7894) );
  MUX2X1 U9813 ( .B(n7898), .A(n7899), .S(n8506), .Y(n7897) );
  MUX2X1 U9814 ( .B(n7901), .A(n7902), .S(n8506), .Y(n7900) );
  MUX2X1 U9815 ( .B(n7904), .A(n7905), .S(n8506), .Y(n7903) );
  MUX2X1 U9816 ( .B(n7907), .A(n7908), .S(n8506), .Y(n7906) );
  MUX2X1 U9817 ( .B(n7910), .A(n7911), .S(N16), .Y(n7909) );
  MUX2X1 U9818 ( .B(n7913), .A(n7914), .S(n8506), .Y(n7912) );
  MUX2X1 U9819 ( .B(n7916), .A(n7917), .S(n8506), .Y(n7915) );
  MUX2X1 U9820 ( .B(n7919), .A(n7920), .S(n8506), .Y(n7918) );
  MUX2X1 U9821 ( .B(n7922), .A(n7923), .S(n8506), .Y(n7921) );
  MUX2X1 U9822 ( .B(n7925), .A(n7926), .S(N16), .Y(n7924) );
  MUX2X1 U9823 ( .B(n7928), .A(n7929), .S(n8507), .Y(n7927) );
  MUX2X1 U9824 ( .B(n7931), .A(n7932), .S(n8507), .Y(n7930) );
  MUX2X1 U9825 ( .B(n7934), .A(n7935), .S(n8507), .Y(n7933) );
  MUX2X1 U9826 ( .B(n7937), .A(n7938), .S(n8507), .Y(n7936) );
  MUX2X1 U9827 ( .B(n7940), .A(n7941), .S(N16), .Y(n7939) );
  MUX2X1 U9828 ( .B(n7943), .A(n7944), .S(n8507), .Y(n7942) );
  MUX2X1 U9829 ( .B(n7946), .A(n7947), .S(n8507), .Y(n7945) );
  MUX2X1 U9830 ( .B(n7949), .A(n7950), .S(n8507), .Y(n7948) );
  MUX2X1 U9831 ( .B(n7952), .A(n7953), .S(n8507), .Y(n7951) );
  MUX2X1 U9832 ( .B(n7955), .A(n7956), .S(N16), .Y(n7954) );
  MUX2X1 U9833 ( .B(n7958), .A(n7959), .S(n8507), .Y(n7957) );
  MUX2X1 U9834 ( .B(n7961), .A(n7962), .S(n8507), .Y(n7960) );
  MUX2X1 U9835 ( .B(n7964), .A(n7965), .S(n8507), .Y(n7963) );
  MUX2X1 U9836 ( .B(n7967), .A(n7968), .S(n8507), .Y(n7966) );
  MUX2X1 U9837 ( .B(n7970), .A(n7971), .S(N16), .Y(n7969) );
  MUX2X1 U9838 ( .B(n7973), .A(n7974), .S(n8508), .Y(n7972) );
  MUX2X1 U9839 ( .B(n7976), .A(n7977), .S(n8508), .Y(n7975) );
  MUX2X1 U9840 ( .B(n7979), .A(n7980), .S(n8508), .Y(n7978) );
  MUX2X1 U9841 ( .B(n7982), .A(n7983), .S(n8508), .Y(n7981) );
  MUX2X1 U9842 ( .B(n7985), .A(n7986), .S(N16), .Y(n7984) );
  MUX2X1 U9843 ( .B(n7988), .A(n7989), .S(n8508), .Y(n7987) );
  MUX2X1 U9844 ( .B(n7991), .A(n7992), .S(n8508), .Y(n7990) );
  MUX2X1 U9845 ( .B(n7994), .A(n7995), .S(n8508), .Y(n7993) );
  MUX2X1 U9846 ( .B(n7997), .A(n7998), .S(n8508), .Y(n7996) );
  MUX2X1 U9847 ( .B(n8000), .A(n8001), .S(N16), .Y(n7999) );
  MUX2X1 U9848 ( .B(n8003), .A(n8004), .S(n8508), .Y(n8002) );
  MUX2X1 U9849 ( .B(n8006), .A(n8007), .S(n8508), .Y(n8005) );
  MUX2X1 U9850 ( .B(n8009), .A(n8010), .S(n8508), .Y(n8008) );
  MUX2X1 U9851 ( .B(n8012), .A(n8013), .S(n8508), .Y(n8011) );
  MUX2X1 U9852 ( .B(n8015), .A(n8016), .S(N16), .Y(n8014) );
  MUX2X1 U9853 ( .B(n8018), .A(n8019), .S(n8509), .Y(n8017) );
  MUX2X1 U9854 ( .B(n8021), .A(n8022), .S(n8509), .Y(n8020) );
  MUX2X1 U9855 ( .B(n8024), .A(n8025), .S(n8509), .Y(n8023) );
  MUX2X1 U9856 ( .B(n8027), .A(n8028), .S(n8509), .Y(n8026) );
  MUX2X1 U9857 ( .B(n8030), .A(n8031), .S(N16), .Y(n8029) );
  MUX2X1 U9858 ( .B(n8033), .A(n8034), .S(n8509), .Y(n8032) );
  MUX2X1 U9859 ( .B(n8036), .A(n8037), .S(n8509), .Y(n8035) );
  MUX2X1 U9860 ( .B(n8039), .A(n8040), .S(n8509), .Y(n8038) );
  MUX2X1 U9861 ( .B(n8042), .A(n8043), .S(n8509), .Y(n8041) );
  MUX2X1 U9862 ( .B(n8045), .A(n8046), .S(N16), .Y(n8044) );
  MUX2X1 U9863 ( .B(n8048), .A(n8049), .S(n8509), .Y(n8047) );
  MUX2X1 U9864 ( .B(n8051), .A(n8052), .S(n8509), .Y(n8050) );
  MUX2X1 U9865 ( .B(n8054), .A(n8055), .S(n8509), .Y(n8053) );
  MUX2X1 U9866 ( .B(n8057), .A(n8058), .S(n8509), .Y(n8056) );
  MUX2X1 U9867 ( .B(n8060), .A(n8061), .S(N16), .Y(n8059) );
  MUX2X1 U9868 ( .B(n8063), .A(n8064), .S(n8510), .Y(n8062) );
  MUX2X1 U9869 ( .B(n8066), .A(n8067), .S(n8510), .Y(n8065) );
  MUX2X1 U9870 ( .B(n8069), .A(n8070), .S(n8510), .Y(n8068) );
  MUX2X1 U9871 ( .B(n8072), .A(n8073), .S(n8510), .Y(n8071) );
  MUX2X1 U9872 ( .B(n8075), .A(n8076), .S(N16), .Y(n8074) );
  MUX2X1 U9873 ( .B(n8078), .A(n8079), .S(n8510), .Y(n8077) );
  MUX2X1 U9874 ( .B(n8081), .A(n8082), .S(n8510), .Y(n8080) );
  MUX2X1 U9875 ( .B(n8084), .A(n8085), .S(n8510), .Y(n8083) );
  MUX2X1 U9876 ( .B(n8087), .A(n8088), .S(n8510), .Y(n8086) );
  MUX2X1 U9877 ( .B(n8090), .A(n8091), .S(N16), .Y(n8089) );
  MUX2X1 U9878 ( .B(n8093), .A(n8094), .S(n8510), .Y(n8092) );
  MUX2X1 U9879 ( .B(n8096), .A(n8097), .S(n8510), .Y(n8095) );
  MUX2X1 U9880 ( .B(n8099), .A(n8100), .S(n8510), .Y(n8098) );
  MUX2X1 U9881 ( .B(n8102), .A(n8103), .S(n8510), .Y(n8101) );
  MUX2X1 U9882 ( .B(n8105), .A(n8106), .S(N16), .Y(n8104) );
  MUX2X1 U9883 ( .B(n8108), .A(n8109), .S(n8511), .Y(n8107) );
  MUX2X1 U9884 ( .B(n8111), .A(n8112), .S(n8511), .Y(n8110) );
  MUX2X1 U9885 ( .B(n8114), .A(n8115), .S(n8511), .Y(n8113) );
  MUX2X1 U9886 ( .B(n8117), .A(n8118), .S(n8511), .Y(n8116) );
  MUX2X1 U9887 ( .B(n8120), .A(n8121), .S(N16), .Y(n8119) );
  MUX2X1 U9888 ( .B(n8123), .A(n8124), .S(n8511), .Y(n8122) );
  MUX2X1 U9889 ( .B(n8126), .A(n8127), .S(n8511), .Y(n8125) );
  MUX2X1 U9890 ( .B(n8129), .A(n8130), .S(n8511), .Y(n8128) );
  MUX2X1 U9891 ( .B(n8132), .A(n8133), .S(n8511), .Y(n8131) );
  MUX2X1 U9892 ( .B(n8135), .A(n8136), .S(N16), .Y(n8134) );
  MUX2X1 U9893 ( .B(n8138), .A(n8139), .S(n8511), .Y(n8137) );
  MUX2X1 U9894 ( .B(n8141), .A(n8142), .S(n8511), .Y(n8140) );
  MUX2X1 U9895 ( .B(n8144), .A(n8145), .S(n8511), .Y(n8143) );
  MUX2X1 U9896 ( .B(n8147), .A(n8148), .S(n8511), .Y(n8146) );
  MUX2X1 U9897 ( .B(n8150), .A(n8151), .S(N16), .Y(n8149) );
  MUX2X1 U9898 ( .B(n8153), .A(n8154), .S(n8512), .Y(n8152) );
  MUX2X1 U9899 ( .B(n8156), .A(n8157), .S(n8512), .Y(n8155) );
  MUX2X1 U9900 ( .B(n8159), .A(n8160), .S(n8512), .Y(n8158) );
  MUX2X1 U9901 ( .B(n8162), .A(n8163), .S(n8512), .Y(n8161) );
  MUX2X1 U9902 ( .B(n8165), .A(n8166), .S(N16), .Y(n8164) );
  MUX2X1 U9903 ( .B(n8168), .A(n8169), .S(n8512), .Y(n8167) );
  MUX2X1 U9904 ( .B(n8171), .A(n8172), .S(n8512), .Y(n8170) );
  MUX2X1 U9905 ( .B(n8174), .A(n8175), .S(n8512), .Y(n8173) );
  MUX2X1 U9906 ( .B(n8177), .A(n8178), .S(n8512), .Y(n8176) );
  MUX2X1 U9907 ( .B(n8180), .A(n8181), .S(N16), .Y(n8179) );
  MUX2X1 U9908 ( .B(n8183), .A(n8184), .S(n8512), .Y(n8182) );
  MUX2X1 U9909 ( .B(n8186), .A(n8187), .S(n8512), .Y(n8185) );
  MUX2X1 U9910 ( .B(n8189), .A(n8190), .S(n8512), .Y(n8188) );
  MUX2X1 U9911 ( .B(n8192), .A(n8193), .S(n8512), .Y(n8191) );
  MUX2X1 U9912 ( .B(n8195), .A(n8196), .S(N16), .Y(n8194) );
  MUX2X1 U9913 ( .B(n8198), .A(n8199), .S(n8513), .Y(n8197) );
  MUX2X1 U9914 ( .B(n8201), .A(n8202), .S(n8513), .Y(n8200) );
  MUX2X1 U9915 ( .B(n8204), .A(n8205), .S(n8513), .Y(n8203) );
  MUX2X1 U9916 ( .B(n8207), .A(n8208), .S(n8513), .Y(n8206) );
  MUX2X1 U9917 ( .B(n8210), .A(n8211), .S(N16), .Y(n8209) );
  MUX2X1 U9918 ( .B(n8213), .A(n8214), .S(n8513), .Y(n8212) );
  MUX2X1 U9919 ( .B(n8216), .A(n8217), .S(n8513), .Y(n8215) );
  MUX2X1 U9920 ( .B(n8219), .A(n8220), .S(n8513), .Y(n8218) );
  MUX2X1 U9921 ( .B(n8222), .A(n8223), .S(n8513), .Y(n8221) );
  MUX2X1 U9922 ( .B(n8225), .A(n8226), .S(N16), .Y(n8224) );
  MUX2X1 U9923 ( .B(n8228), .A(n8229), .S(n8513), .Y(n8227) );
  MUX2X1 U9924 ( .B(n8231), .A(n8232), .S(n8513), .Y(n8230) );
  MUX2X1 U9925 ( .B(n8234), .A(n8235), .S(n8513), .Y(n8233) );
  MUX2X1 U9926 ( .B(n8237), .A(n8238), .S(n8513), .Y(n8236) );
  MUX2X1 U9927 ( .B(n8240), .A(n8241), .S(N16), .Y(n8239) );
  MUX2X1 U9928 ( .B(n8243), .A(n8244), .S(n8514), .Y(n8242) );
  MUX2X1 U9929 ( .B(n8246), .A(n8247), .S(n8514), .Y(n8245) );
  MUX2X1 U9930 ( .B(n8249), .A(n8250), .S(n8514), .Y(n8248) );
  MUX2X1 U9931 ( .B(n8252), .A(n8253), .S(n8514), .Y(n8251) );
  MUX2X1 U9932 ( .B(n8255), .A(n8256), .S(N16), .Y(n8254) );
  MUX2X1 U9933 ( .B(n8258), .A(n8259), .S(n8514), .Y(n8257) );
  MUX2X1 U9934 ( .B(n8261), .A(n8262), .S(n8514), .Y(n8260) );
  MUX2X1 U9935 ( .B(n8264), .A(n8265), .S(n8514), .Y(n8263) );
  MUX2X1 U9936 ( .B(n8267), .A(n8268), .S(n8514), .Y(n8266) );
  MUX2X1 U9937 ( .B(n8270), .A(n8271), .S(N16), .Y(n8269) );
  MUX2X1 U9938 ( .B(n8273), .A(n8274), .S(n8514), .Y(n8272) );
  MUX2X1 U9939 ( .B(n8276), .A(n8277), .S(n8514), .Y(n8275) );
  MUX2X1 U9940 ( .B(n8279), .A(n8280), .S(n8514), .Y(n8278) );
  MUX2X1 U9941 ( .B(n8282), .A(n8283), .S(n8514), .Y(n8281) );
  MUX2X1 U9942 ( .B(n8285), .A(n8286), .S(N16), .Y(n8284) );
  MUX2X1 U9943 ( .B(\RF[30][0] ), .A(\RF[31][0] ), .S(n8371), .Y(n6369) );
  MUX2X1 U9944 ( .B(\RF[28][0] ), .A(\RF[29][0] ), .S(n8371), .Y(n6368) );
  MUX2X1 U9945 ( .B(\RF[26][0] ), .A(\RF[27][0] ), .S(n8371), .Y(n6372) );
  MUX2X1 U9946 ( .B(\RF[24][0] ), .A(\RF[25][0] ), .S(n8371), .Y(n6371) );
  MUX2X1 U9947 ( .B(n6370), .A(n6367), .S(N15), .Y(n6381) );
  MUX2X1 U9948 ( .B(\RF[22][0] ), .A(\RF[23][0] ), .S(n8372), .Y(n6375) );
  MUX2X1 U9949 ( .B(\RF[20][0] ), .A(\RF[21][0] ), .S(n8372), .Y(n6374) );
  MUX2X1 U9950 ( .B(\RF[18][0] ), .A(\RF[19][0] ), .S(n8372), .Y(n6378) );
  MUX2X1 U9951 ( .B(\RF[16][0] ), .A(\RF[17][0] ), .S(n8372), .Y(n6377) );
  MUX2X1 U9952 ( .B(n6376), .A(n6373), .S(N15), .Y(n6380) );
  MUX2X1 U9953 ( .B(\RF[14][0] ), .A(\RF[15][0] ), .S(n8372), .Y(n6384) );
  MUX2X1 U9954 ( .B(\RF[12][0] ), .A(\RF[13][0] ), .S(n8372), .Y(n6383) );
  MUX2X1 U9955 ( .B(\RF[10][0] ), .A(\RF[11][0] ), .S(n8372), .Y(n6387) );
  MUX2X1 U9956 ( .B(\RF[8][0] ), .A(\RF[9][0] ), .S(n8372), .Y(n6386) );
  MUX2X1 U9957 ( .B(n6385), .A(n6382), .S(N15), .Y(n6396) );
  MUX2X1 U9958 ( .B(\RF[6][0] ), .A(\RF[7][0] ), .S(n8372), .Y(n6390) );
  MUX2X1 U9959 ( .B(\RF[4][0] ), .A(\RF[5][0] ), .S(n8372), .Y(n6389) );
  MUX2X1 U9960 ( .B(\RF[2][0] ), .A(\RF[3][0] ), .S(n8372), .Y(n6393) );
  MUX2X1 U9961 ( .B(\RF[0][0] ), .A(\RF[1][0] ), .S(n8372), .Y(n6392) );
  MUX2X1 U9962 ( .B(n6391), .A(n6388), .S(N15), .Y(n6395) );
  MUX2X1 U9963 ( .B(n6394), .A(n6379), .S(N17), .Y(n8287) );
  MUX2X1 U9964 ( .B(\RF[30][1] ), .A(\RF[31][1] ), .S(n8373), .Y(n6399) );
  MUX2X1 U9965 ( .B(\RF[28][1] ), .A(\RF[29][1] ), .S(n8373), .Y(n6398) );
  MUX2X1 U9966 ( .B(\RF[26][1] ), .A(\RF[27][1] ), .S(n8373), .Y(n6402) );
  MUX2X1 U9967 ( .B(\RF[24][1] ), .A(\RF[25][1] ), .S(n8373), .Y(n6401) );
  MUX2X1 U9968 ( .B(n6400), .A(n6397), .S(n8517), .Y(n6411) );
  MUX2X1 U9969 ( .B(\RF[22][1] ), .A(\RF[23][1] ), .S(n8373), .Y(n6405) );
  MUX2X1 U9970 ( .B(\RF[20][1] ), .A(\RF[21][1] ), .S(n8373), .Y(n6404) );
  MUX2X1 U9971 ( .B(\RF[18][1] ), .A(\RF[19][1] ), .S(n8373), .Y(n6408) );
  MUX2X1 U9972 ( .B(\RF[16][1] ), .A(\RF[17][1] ), .S(n8373), .Y(n6407) );
  MUX2X1 U9973 ( .B(n6406), .A(n6403), .S(n8517), .Y(n6410) );
  MUX2X1 U9974 ( .B(\RF[14][1] ), .A(\RF[15][1] ), .S(n8373), .Y(n6414) );
  MUX2X1 U9975 ( .B(\RF[12][1] ), .A(\RF[13][1] ), .S(n8373), .Y(n6413) );
  MUX2X1 U9976 ( .B(\RF[10][1] ), .A(\RF[11][1] ), .S(n8373), .Y(n6417) );
  MUX2X1 U9977 ( .B(\RF[8][1] ), .A(\RF[9][1] ), .S(n8373), .Y(n6416) );
  MUX2X1 U9978 ( .B(n6415), .A(n6412), .S(n8517), .Y(n6426) );
  MUX2X1 U9979 ( .B(\RF[6][1] ), .A(\RF[7][1] ), .S(n8374), .Y(n6420) );
  MUX2X1 U9980 ( .B(\RF[4][1] ), .A(\RF[5][1] ), .S(n8374), .Y(n6419) );
  MUX2X1 U9981 ( .B(\RF[2][1] ), .A(\RF[3][1] ), .S(n8374), .Y(n6423) );
  MUX2X1 U9982 ( .B(\RF[0][1] ), .A(\RF[1][1] ), .S(n8374), .Y(n6422) );
  MUX2X1 U9983 ( .B(n6421), .A(n6418), .S(n8517), .Y(n6425) );
  MUX2X1 U9984 ( .B(n6424), .A(n6409), .S(N17), .Y(n8288) );
  MUX2X1 U9985 ( .B(\RF[30][2] ), .A(\RF[31][2] ), .S(n8374), .Y(n6429) );
  MUX2X1 U9986 ( .B(\RF[28][2] ), .A(\RF[29][2] ), .S(n8374), .Y(n6428) );
  MUX2X1 U9987 ( .B(\RF[26][2] ), .A(\RF[27][2] ), .S(n8374), .Y(n6432) );
  MUX2X1 U9988 ( .B(\RF[24][2] ), .A(\RF[25][2] ), .S(n8374), .Y(n6431) );
  MUX2X1 U9989 ( .B(n6430), .A(n6427), .S(n8517), .Y(n6441) );
  MUX2X1 U9990 ( .B(\RF[22][2] ), .A(\RF[23][2] ), .S(n8374), .Y(n6435) );
  MUX2X1 U9991 ( .B(\RF[20][2] ), .A(\RF[21][2] ), .S(n8374), .Y(n6434) );
  MUX2X1 U9992 ( .B(\RF[18][2] ), .A(\RF[19][2] ), .S(n8374), .Y(n6438) );
  MUX2X1 U9993 ( .B(\RF[16][2] ), .A(\RF[17][2] ), .S(n8374), .Y(n6437) );
  MUX2X1 U9994 ( .B(n6436), .A(n6433), .S(n8517), .Y(n6440) );
  MUX2X1 U9995 ( .B(\RF[14][2] ), .A(\RF[15][2] ), .S(n8375), .Y(n6444) );
  MUX2X1 U9996 ( .B(\RF[12][2] ), .A(\RF[13][2] ), .S(n8375), .Y(n6443) );
  MUX2X1 U9997 ( .B(\RF[10][2] ), .A(\RF[11][2] ), .S(n8375), .Y(n6447) );
  MUX2X1 U9998 ( .B(\RF[8][2] ), .A(\RF[9][2] ), .S(n8375), .Y(n6446) );
  MUX2X1 U9999 ( .B(n6445), .A(n6442), .S(n8517), .Y(n6456) );
  MUX2X1 U10000 ( .B(\RF[6][2] ), .A(\RF[7][2] ), .S(n8375), .Y(n6450) );
  MUX2X1 U10001 ( .B(\RF[4][2] ), .A(\RF[5][2] ), .S(n8375), .Y(n6449) );
  MUX2X1 U10002 ( .B(\RF[2][2] ), .A(\RF[3][2] ), .S(n8375), .Y(n6453) );
  MUX2X1 U10003 ( .B(\RF[0][2] ), .A(\RF[1][2] ), .S(n8375), .Y(n6452) );
  MUX2X1 U10004 ( .B(n6451), .A(n6448), .S(n8517), .Y(n6455) );
  MUX2X1 U10005 ( .B(n6454), .A(n6439), .S(N17), .Y(n8289) );
  MUX2X1 U10006 ( .B(\RF[30][3] ), .A(\RF[31][3] ), .S(n8375), .Y(n6459) );
  MUX2X1 U10007 ( .B(\RF[28][3] ), .A(\RF[29][3] ), .S(n8375), .Y(n6458) );
  MUX2X1 U10008 ( .B(\RF[26][3] ), .A(\RF[27][3] ), .S(n8375), .Y(n6462) );
  MUX2X1 U10009 ( .B(\RF[24][3] ), .A(\RF[25][3] ), .S(n8375), .Y(n6461) );
  MUX2X1 U10010 ( .B(n6460), .A(n6457), .S(n8517), .Y(n6471) );
  MUX2X1 U10011 ( .B(\RF[22][3] ), .A(\RF[23][3] ), .S(n8376), .Y(n6465) );
  MUX2X1 U10012 ( .B(\RF[20][3] ), .A(\RF[21][3] ), .S(n8376), .Y(n6464) );
  MUX2X1 U10013 ( .B(\RF[18][3] ), .A(\RF[19][3] ), .S(n8376), .Y(n6468) );
  MUX2X1 U10014 ( .B(\RF[16][3] ), .A(\RF[17][3] ), .S(n8376), .Y(n6467) );
  MUX2X1 U10015 ( .B(n6466), .A(n6463), .S(n8517), .Y(n6470) );
  MUX2X1 U10016 ( .B(\RF[14][3] ), .A(\RF[15][3] ), .S(n8376), .Y(n6474) );
  MUX2X1 U10017 ( .B(\RF[12][3] ), .A(\RF[13][3] ), .S(n8376), .Y(n6473) );
  MUX2X1 U10018 ( .B(\RF[10][3] ), .A(\RF[11][3] ), .S(n8376), .Y(n6477) );
  MUX2X1 U10019 ( .B(\RF[8][3] ), .A(\RF[9][3] ), .S(n8376), .Y(n6476) );
  MUX2X1 U10020 ( .B(n6475), .A(n6472), .S(n8517), .Y(n6486) );
  MUX2X1 U10021 ( .B(\RF[6][3] ), .A(\RF[7][3] ), .S(n8376), .Y(n6480) );
  MUX2X1 U10022 ( .B(\RF[4][3] ), .A(\RF[5][3] ), .S(n8376), .Y(n6479) );
  MUX2X1 U10023 ( .B(\RF[2][3] ), .A(\RF[3][3] ), .S(n8376), .Y(n6483) );
  MUX2X1 U10024 ( .B(\RF[0][3] ), .A(\RF[1][3] ), .S(n8376), .Y(n6482) );
  MUX2X1 U10025 ( .B(n6481), .A(n6478), .S(n8517), .Y(n6485) );
  MUX2X1 U10026 ( .B(n6484), .A(n6469), .S(N17), .Y(n8290) );
  MUX2X1 U10027 ( .B(\RF[30][4] ), .A(\RF[31][4] ), .S(n8377), .Y(n6489) );
  MUX2X1 U10028 ( .B(\RF[28][4] ), .A(\RF[29][4] ), .S(n8377), .Y(n6488) );
  MUX2X1 U10029 ( .B(\RF[26][4] ), .A(\RF[27][4] ), .S(n8377), .Y(n6492) );
  MUX2X1 U10030 ( .B(\RF[24][4] ), .A(\RF[25][4] ), .S(n8377), .Y(n6491) );
  MUX2X1 U10031 ( .B(n6490), .A(n6487), .S(n8518), .Y(n6501) );
  MUX2X1 U10032 ( .B(\RF[22][4] ), .A(\RF[23][4] ), .S(n8377), .Y(n6495) );
  MUX2X1 U10033 ( .B(\RF[20][4] ), .A(\RF[21][4] ), .S(n8377), .Y(n6494) );
  MUX2X1 U10034 ( .B(\RF[18][4] ), .A(\RF[19][4] ), .S(n8377), .Y(n6498) );
  MUX2X1 U10035 ( .B(\RF[16][4] ), .A(\RF[17][4] ), .S(n8377), .Y(n6497) );
  MUX2X1 U10036 ( .B(n6496), .A(n6493), .S(n8518), .Y(n6500) );
  MUX2X1 U10037 ( .B(\RF[14][4] ), .A(\RF[15][4] ), .S(n8377), .Y(n6504) );
  MUX2X1 U10038 ( .B(\RF[12][4] ), .A(\RF[13][4] ), .S(n8377), .Y(n6503) );
  MUX2X1 U10039 ( .B(\RF[10][4] ), .A(\RF[11][4] ), .S(n8377), .Y(n6507) );
  MUX2X1 U10040 ( .B(\RF[8][4] ), .A(\RF[9][4] ), .S(n8377), .Y(n6506) );
  MUX2X1 U10041 ( .B(n6505), .A(n6502), .S(n8518), .Y(n6516) );
  MUX2X1 U10042 ( .B(\RF[6][4] ), .A(\RF[7][4] ), .S(n8378), .Y(n6510) );
  MUX2X1 U10043 ( .B(\RF[4][4] ), .A(\RF[5][4] ), .S(n8378), .Y(n6509) );
  MUX2X1 U10044 ( .B(\RF[2][4] ), .A(\RF[3][4] ), .S(n8378), .Y(n6513) );
  MUX2X1 U10045 ( .B(\RF[0][4] ), .A(\RF[1][4] ), .S(n8378), .Y(n6512) );
  MUX2X1 U10046 ( .B(n6511), .A(n6508), .S(n8518), .Y(n6515) );
  MUX2X1 U10047 ( .B(n6514), .A(n6499), .S(N17), .Y(n8291) );
  MUX2X1 U10048 ( .B(\RF[30][5] ), .A(\RF[31][5] ), .S(n8378), .Y(n6519) );
  MUX2X1 U10049 ( .B(\RF[28][5] ), .A(\RF[29][5] ), .S(n8378), .Y(n6518) );
  MUX2X1 U10050 ( .B(\RF[26][5] ), .A(\RF[27][5] ), .S(n8378), .Y(n6522) );
  MUX2X1 U10051 ( .B(\RF[24][5] ), .A(\RF[25][5] ), .S(n8378), .Y(n6521) );
  MUX2X1 U10052 ( .B(n6520), .A(n6517), .S(n8518), .Y(n6531) );
  MUX2X1 U10053 ( .B(\RF[22][5] ), .A(\RF[23][5] ), .S(n8378), .Y(n6525) );
  MUX2X1 U10054 ( .B(\RF[20][5] ), .A(\RF[21][5] ), .S(n8378), .Y(n6524) );
  MUX2X1 U10055 ( .B(\RF[18][5] ), .A(\RF[19][5] ), .S(n8378), .Y(n6528) );
  MUX2X1 U10056 ( .B(\RF[16][5] ), .A(\RF[17][5] ), .S(n8378), .Y(n6527) );
  MUX2X1 U10057 ( .B(n6526), .A(n6523), .S(n8518), .Y(n6530) );
  MUX2X1 U10058 ( .B(\RF[14][5] ), .A(\RF[15][5] ), .S(n8379), .Y(n6534) );
  MUX2X1 U10059 ( .B(\RF[12][5] ), .A(\RF[13][5] ), .S(n8379), .Y(n6533) );
  MUX2X1 U10060 ( .B(\RF[10][5] ), .A(\RF[11][5] ), .S(n8379), .Y(n6537) );
  MUX2X1 U10061 ( .B(\RF[8][5] ), .A(\RF[9][5] ), .S(n8379), .Y(n6536) );
  MUX2X1 U10062 ( .B(n6535), .A(n6532), .S(n8518), .Y(n6546) );
  MUX2X1 U10063 ( .B(\RF[6][5] ), .A(\RF[7][5] ), .S(n8379), .Y(n6540) );
  MUX2X1 U10064 ( .B(\RF[4][5] ), .A(\RF[5][5] ), .S(n8379), .Y(n6539) );
  MUX2X1 U10065 ( .B(\RF[2][5] ), .A(\RF[3][5] ), .S(n8379), .Y(n6543) );
  MUX2X1 U10066 ( .B(\RF[0][5] ), .A(\RF[1][5] ), .S(n8379), .Y(n6542) );
  MUX2X1 U10067 ( .B(n6541), .A(n6538), .S(n8518), .Y(n6545) );
  MUX2X1 U10068 ( .B(n6544), .A(n6529), .S(N17), .Y(n8292) );
  MUX2X1 U10069 ( .B(\RF[30][6] ), .A(\RF[31][6] ), .S(n8379), .Y(n6549) );
  MUX2X1 U10070 ( .B(\RF[28][6] ), .A(\RF[29][6] ), .S(n8379), .Y(n6548) );
  MUX2X1 U10071 ( .B(\RF[26][6] ), .A(\RF[27][6] ), .S(n8379), .Y(n6552) );
  MUX2X1 U10072 ( .B(\RF[24][6] ), .A(\RF[25][6] ), .S(n8379), .Y(n6551) );
  MUX2X1 U10073 ( .B(n6550), .A(n6547), .S(n8518), .Y(n6561) );
  MUX2X1 U10074 ( .B(\RF[22][6] ), .A(\RF[23][6] ), .S(n8380), .Y(n6555) );
  MUX2X1 U10075 ( .B(\RF[20][6] ), .A(\RF[21][6] ), .S(n8380), .Y(n6554) );
  MUX2X1 U10076 ( .B(\RF[18][6] ), .A(\RF[19][6] ), .S(n8380), .Y(n6558) );
  MUX2X1 U10077 ( .B(\RF[16][6] ), .A(\RF[17][6] ), .S(n8380), .Y(n6557) );
  MUX2X1 U10078 ( .B(n6556), .A(n6553), .S(n8518), .Y(n6560) );
  MUX2X1 U10079 ( .B(\RF[14][6] ), .A(\RF[15][6] ), .S(n8380), .Y(n6564) );
  MUX2X1 U10080 ( .B(\RF[12][6] ), .A(\RF[13][6] ), .S(n8380), .Y(n6563) );
  MUX2X1 U10081 ( .B(\RF[10][6] ), .A(\RF[11][6] ), .S(n8380), .Y(n6567) );
  MUX2X1 U10082 ( .B(\RF[8][6] ), .A(\RF[9][6] ), .S(n8380), .Y(n6566) );
  MUX2X1 U10083 ( .B(n6565), .A(n6562), .S(n8518), .Y(n6576) );
  MUX2X1 U10084 ( .B(\RF[6][6] ), .A(\RF[7][6] ), .S(n8380), .Y(n6570) );
  MUX2X1 U10085 ( .B(\RF[4][6] ), .A(\RF[5][6] ), .S(n8380), .Y(n6569) );
  MUX2X1 U10086 ( .B(\RF[2][6] ), .A(\RF[3][6] ), .S(n8380), .Y(n6573) );
  MUX2X1 U10087 ( .B(\RF[0][6] ), .A(\RF[1][6] ), .S(n8380), .Y(n6572) );
  MUX2X1 U10088 ( .B(n6571), .A(n6568), .S(n8518), .Y(n6575) );
  MUX2X1 U10089 ( .B(n6574), .A(n6559), .S(N17), .Y(n8293) );
  MUX2X1 U10090 ( .B(\RF[30][7] ), .A(\RF[31][7] ), .S(n8381), .Y(n6579) );
  MUX2X1 U10091 ( .B(\RF[28][7] ), .A(\RF[29][7] ), .S(n8381), .Y(n6578) );
  MUX2X1 U10092 ( .B(\RF[26][7] ), .A(\RF[27][7] ), .S(n8381), .Y(n6582) );
  MUX2X1 U10093 ( .B(\RF[24][7] ), .A(\RF[25][7] ), .S(n8381), .Y(n6581) );
  MUX2X1 U10094 ( .B(n6580), .A(n6577), .S(n8519), .Y(n6591) );
  MUX2X1 U10095 ( .B(\RF[22][7] ), .A(\RF[23][7] ), .S(n8381), .Y(n6585) );
  MUX2X1 U10096 ( .B(\RF[20][7] ), .A(\RF[21][7] ), .S(n8381), .Y(n6584) );
  MUX2X1 U10097 ( .B(\RF[18][7] ), .A(\RF[19][7] ), .S(n8381), .Y(n6588) );
  MUX2X1 U10098 ( .B(\RF[16][7] ), .A(\RF[17][7] ), .S(n8381), .Y(n6587) );
  MUX2X1 U10099 ( .B(n6586), .A(n6583), .S(n8519), .Y(n6590) );
  MUX2X1 U10100 ( .B(\RF[14][7] ), .A(\RF[15][7] ), .S(n8381), .Y(n6594) );
  MUX2X1 U10101 ( .B(\RF[12][7] ), .A(\RF[13][7] ), .S(n8381), .Y(n6593) );
  MUX2X1 U10102 ( .B(\RF[10][7] ), .A(\RF[11][7] ), .S(n8381), .Y(n6597) );
  MUX2X1 U10103 ( .B(\RF[8][7] ), .A(\RF[9][7] ), .S(n8381), .Y(n6596) );
  MUX2X1 U10104 ( .B(n6595), .A(n6592), .S(n8519), .Y(n6606) );
  MUX2X1 U10105 ( .B(\RF[6][7] ), .A(\RF[7][7] ), .S(n8382), .Y(n6600) );
  MUX2X1 U10106 ( .B(\RF[4][7] ), .A(\RF[5][7] ), .S(n8382), .Y(n6599) );
  MUX2X1 U10107 ( .B(\RF[2][7] ), .A(\RF[3][7] ), .S(n8382), .Y(n6603) );
  MUX2X1 U10108 ( .B(\RF[0][7] ), .A(\RF[1][7] ), .S(n8382), .Y(n6602) );
  MUX2X1 U10109 ( .B(n6601), .A(n6598), .S(n8519), .Y(n6605) );
  MUX2X1 U10110 ( .B(n6604), .A(n6589), .S(N17), .Y(n8294) );
  MUX2X1 U10111 ( .B(\RF[30][8] ), .A(\RF[31][8] ), .S(n8382), .Y(n6609) );
  MUX2X1 U10112 ( .B(\RF[28][8] ), .A(\RF[29][8] ), .S(n8382), .Y(n6608) );
  MUX2X1 U10113 ( .B(\RF[26][8] ), .A(\RF[27][8] ), .S(n8382), .Y(n6612) );
  MUX2X1 U10114 ( .B(\RF[24][8] ), .A(\RF[25][8] ), .S(n8382), .Y(n6611) );
  MUX2X1 U10115 ( .B(n6610), .A(n6607), .S(n8519), .Y(n6621) );
  MUX2X1 U10116 ( .B(\RF[22][8] ), .A(\RF[23][8] ), .S(n8382), .Y(n6615) );
  MUX2X1 U10117 ( .B(\RF[20][8] ), .A(\RF[21][8] ), .S(n8382), .Y(n6614) );
  MUX2X1 U10118 ( .B(\RF[18][8] ), .A(\RF[19][8] ), .S(n8382), .Y(n6618) );
  MUX2X1 U10119 ( .B(\RF[16][8] ), .A(\RF[17][8] ), .S(n8382), .Y(n6617) );
  MUX2X1 U10120 ( .B(n6616), .A(n6613), .S(n8519), .Y(n6620) );
  MUX2X1 U10121 ( .B(\RF[14][8] ), .A(\RF[15][8] ), .S(n8383), .Y(n6624) );
  MUX2X1 U10122 ( .B(\RF[12][8] ), .A(\RF[13][8] ), .S(n8383), .Y(n6623) );
  MUX2X1 U10123 ( .B(\RF[10][8] ), .A(\RF[11][8] ), .S(n8383), .Y(n6627) );
  MUX2X1 U10124 ( .B(\RF[8][8] ), .A(\RF[9][8] ), .S(n8383), .Y(n6626) );
  MUX2X1 U10125 ( .B(n6625), .A(n6622), .S(n8519), .Y(n6636) );
  MUX2X1 U10126 ( .B(\RF[6][8] ), .A(\RF[7][8] ), .S(n8383), .Y(n6630) );
  MUX2X1 U10127 ( .B(\RF[4][8] ), .A(\RF[5][8] ), .S(n8383), .Y(n6629) );
  MUX2X1 U10128 ( .B(\RF[2][8] ), .A(\RF[3][8] ), .S(n8383), .Y(n6633) );
  MUX2X1 U10129 ( .B(\RF[0][8] ), .A(\RF[1][8] ), .S(n8383), .Y(n6632) );
  MUX2X1 U10130 ( .B(n6631), .A(n6628), .S(n8519), .Y(n6635) );
  MUX2X1 U10131 ( .B(n6634), .A(n6619), .S(N17), .Y(n8295) );
  MUX2X1 U10132 ( .B(\RF[30][9] ), .A(\RF[31][9] ), .S(n8383), .Y(n6639) );
  MUX2X1 U10133 ( .B(\RF[28][9] ), .A(\RF[29][9] ), .S(n8383), .Y(n6638) );
  MUX2X1 U10134 ( .B(\RF[26][9] ), .A(\RF[27][9] ), .S(n8383), .Y(n6642) );
  MUX2X1 U10135 ( .B(\RF[24][9] ), .A(\RF[25][9] ), .S(n8383), .Y(n6641) );
  MUX2X1 U10136 ( .B(n6640), .A(n6637), .S(n8519), .Y(n6651) );
  MUX2X1 U10137 ( .B(\RF[22][9] ), .A(\RF[23][9] ), .S(n8384), .Y(n6645) );
  MUX2X1 U10138 ( .B(\RF[20][9] ), .A(\RF[21][9] ), .S(n8384), .Y(n6644) );
  MUX2X1 U10139 ( .B(\RF[18][9] ), .A(\RF[19][9] ), .S(n8384), .Y(n6648) );
  MUX2X1 U10140 ( .B(\RF[16][9] ), .A(\RF[17][9] ), .S(n8384), .Y(n6647) );
  MUX2X1 U10141 ( .B(n6646), .A(n6643), .S(n8519), .Y(n6650) );
  MUX2X1 U10142 ( .B(\RF[14][9] ), .A(\RF[15][9] ), .S(n8384), .Y(n6654) );
  MUX2X1 U10143 ( .B(\RF[12][9] ), .A(\RF[13][9] ), .S(n8384), .Y(n6653) );
  MUX2X1 U10144 ( .B(\RF[10][9] ), .A(\RF[11][9] ), .S(n8384), .Y(n6657) );
  MUX2X1 U10145 ( .B(\RF[8][9] ), .A(\RF[9][9] ), .S(n8384), .Y(n6656) );
  MUX2X1 U10146 ( .B(n6655), .A(n6652), .S(n8519), .Y(n6666) );
  MUX2X1 U10147 ( .B(\RF[6][9] ), .A(\RF[7][9] ), .S(n8384), .Y(n6660) );
  MUX2X1 U10148 ( .B(\RF[4][9] ), .A(\RF[5][9] ), .S(n8384), .Y(n6659) );
  MUX2X1 U10149 ( .B(\RF[2][9] ), .A(\RF[3][9] ), .S(n8384), .Y(n6663) );
  MUX2X1 U10150 ( .B(\RF[0][9] ), .A(\RF[1][9] ), .S(n8384), .Y(n6662) );
  MUX2X1 U10151 ( .B(n6661), .A(n6658), .S(n8519), .Y(n6665) );
  MUX2X1 U10152 ( .B(n6664), .A(n6649), .S(N17), .Y(n8296) );
  MUX2X1 U10153 ( .B(\RF[30][10] ), .A(\RF[31][10] ), .S(n8385), .Y(n6669) );
  MUX2X1 U10154 ( .B(\RF[28][10] ), .A(\RF[29][10] ), .S(n8385), .Y(n6668) );
  MUX2X1 U10155 ( .B(\RF[26][10] ), .A(\RF[27][10] ), .S(n8385), .Y(n6672) );
  MUX2X1 U10156 ( .B(\RF[24][10] ), .A(\RF[25][10] ), .S(n8385), .Y(n6671) );
  MUX2X1 U10157 ( .B(n6670), .A(n6667), .S(n8520), .Y(n6681) );
  MUX2X1 U10158 ( .B(\RF[22][10] ), .A(\RF[23][10] ), .S(n8385), .Y(n6675) );
  MUX2X1 U10159 ( .B(\RF[20][10] ), .A(\RF[21][10] ), .S(n8385), .Y(n6674) );
  MUX2X1 U10160 ( .B(\RF[18][10] ), .A(\RF[19][10] ), .S(n8385), .Y(n6678) );
  MUX2X1 U10161 ( .B(\RF[16][10] ), .A(\RF[17][10] ), .S(n8385), .Y(n6677) );
  MUX2X1 U10162 ( .B(n6676), .A(n6673), .S(n8520), .Y(n6680) );
  MUX2X1 U10163 ( .B(\RF[14][10] ), .A(\RF[15][10] ), .S(n8385), .Y(n6684) );
  MUX2X1 U10164 ( .B(\RF[12][10] ), .A(\RF[13][10] ), .S(n8385), .Y(n6683) );
  MUX2X1 U10165 ( .B(\RF[10][10] ), .A(\RF[11][10] ), .S(n8385), .Y(n6687) );
  MUX2X1 U10166 ( .B(\RF[8][10] ), .A(\RF[9][10] ), .S(n8385), .Y(n6686) );
  MUX2X1 U10167 ( .B(n6685), .A(n6682), .S(n8520), .Y(n6696) );
  MUX2X1 U10168 ( .B(\RF[6][10] ), .A(\RF[7][10] ), .S(n8386), .Y(n6690) );
  MUX2X1 U10169 ( .B(\RF[4][10] ), .A(\RF[5][10] ), .S(n8386), .Y(n6689) );
  MUX2X1 U10170 ( .B(\RF[2][10] ), .A(\RF[3][10] ), .S(n8386), .Y(n6693) );
  MUX2X1 U10171 ( .B(\RF[0][10] ), .A(\RF[1][10] ), .S(n8386), .Y(n6692) );
  MUX2X1 U10172 ( .B(n6691), .A(n6688), .S(n8520), .Y(n6695) );
  MUX2X1 U10173 ( .B(n6694), .A(n6679), .S(N17), .Y(n8297) );
  MUX2X1 U10174 ( .B(\RF[30][11] ), .A(\RF[31][11] ), .S(n8386), .Y(n6699) );
  MUX2X1 U10175 ( .B(\RF[28][11] ), .A(\RF[29][11] ), .S(n8386), .Y(n6698) );
  MUX2X1 U10176 ( .B(\RF[26][11] ), .A(\RF[27][11] ), .S(n8386), .Y(n6702) );
  MUX2X1 U10177 ( .B(\RF[24][11] ), .A(\RF[25][11] ), .S(n8386), .Y(n6701) );
  MUX2X1 U10178 ( .B(n6700), .A(n6697), .S(n8520), .Y(n6711) );
  MUX2X1 U10179 ( .B(\RF[22][11] ), .A(\RF[23][11] ), .S(n8386), .Y(n6705) );
  MUX2X1 U10180 ( .B(\RF[20][11] ), .A(\RF[21][11] ), .S(n8386), .Y(n6704) );
  MUX2X1 U10181 ( .B(\RF[18][11] ), .A(\RF[19][11] ), .S(n8386), .Y(n6708) );
  MUX2X1 U10182 ( .B(\RF[16][11] ), .A(\RF[17][11] ), .S(n8386), .Y(n6707) );
  MUX2X1 U10183 ( .B(n6706), .A(n6703), .S(n8520), .Y(n6710) );
  MUX2X1 U10184 ( .B(\RF[14][11] ), .A(\RF[15][11] ), .S(n8387), .Y(n6714) );
  MUX2X1 U10185 ( .B(\RF[12][11] ), .A(\RF[13][11] ), .S(n8387), .Y(n6713) );
  MUX2X1 U10186 ( .B(\RF[10][11] ), .A(\RF[11][11] ), .S(n8387), .Y(n6717) );
  MUX2X1 U10187 ( .B(\RF[8][11] ), .A(\RF[9][11] ), .S(n8387), .Y(n6716) );
  MUX2X1 U10188 ( .B(n6715), .A(n6712), .S(n8520), .Y(n6726) );
  MUX2X1 U10189 ( .B(\RF[6][11] ), .A(\RF[7][11] ), .S(n8387), .Y(n6720) );
  MUX2X1 U10190 ( .B(\RF[4][11] ), .A(\RF[5][11] ), .S(n8387), .Y(n6719) );
  MUX2X1 U10191 ( .B(\RF[2][11] ), .A(\RF[3][11] ), .S(n8387), .Y(n6723) );
  MUX2X1 U10192 ( .B(\RF[0][11] ), .A(\RF[1][11] ), .S(n8387), .Y(n6722) );
  MUX2X1 U10193 ( .B(n6721), .A(n6718), .S(n8520), .Y(n6725) );
  MUX2X1 U10194 ( .B(n6724), .A(n6709), .S(N17), .Y(n8298) );
  MUX2X1 U10195 ( .B(\RF[30][12] ), .A(\RF[31][12] ), .S(n8387), .Y(n6729) );
  MUX2X1 U10196 ( .B(\RF[28][12] ), .A(\RF[29][12] ), .S(n8387), .Y(n6728) );
  MUX2X1 U10197 ( .B(\RF[26][12] ), .A(\RF[27][12] ), .S(n8387), .Y(n6732) );
  MUX2X1 U10198 ( .B(\RF[24][12] ), .A(\RF[25][12] ), .S(n8387), .Y(n6731) );
  MUX2X1 U10199 ( .B(n6730), .A(n6727), .S(n8520), .Y(n6741) );
  MUX2X1 U10200 ( .B(\RF[22][12] ), .A(\RF[23][12] ), .S(n8388), .Y(n6735) );
  MUX2X1 U10201 ( .B(\RF[20][12] ), .A(\RF[21][12] ), .S(n8388), .Y(n6734) );
  MUX2X1 U10202 ( .B(\RF[18][12] ), .A(\RF[19][12] ), .S(n8388), .Y(n6738) );
  MUX2X1 U10203 ( .B(\RF[16][12] ), .A(\RF[17][12] ), .S(n8388), .Y(n6737) );
  MUX2X1 U10204 ( .B(n6736), .A(n6733), .S(n8520), .Y(n6740) );
  MUX2X1 U10205 ( .B(\RF[14][12] ), .A(\RF[15][12] ), .S(n8388), .Y(n6744) );
  MUX2X1 U10206 ( .B(\RF[12][12] ), .A(\RF[13][12] ), .S(n8388), .Y(n6743) );
  MUX2X1 U10207 ( .B(\RF[10][12] ), .A(\RF[11][12] ), .S(n8388), .Y(n6747) );
  MUX2X1 U10208 ( .B(\RF[8][12] ), .A(\RF[9][12] ), .S(n8388), .Y(n6746) );
  MUX2X1 U10209 ( .B(n6745), .A(n6742), .S(n8520), .Y(n6756) );
  MUX2X1 U10210 ( .B(\RF[6][12] ), .A(\RF[7][12] ), .S(n8388), .Y(n6750) );
  MUX2X1 U10211 ( .B(\RF[4][12] ), .A(\RF[5][12] ), .S(n8388), .Y(n6749) );
  MUX2X1 U10212 ( .B(\RF[2][12] ), .A(\RF[3][12] ), .S(n8388), .Y(n6753) );
  MUX2X1 U10213 ( .B(\RF[0][12] ), .A(\RF[1][12] ), .S(n8388), .Y(n6752) );
  MUX2X1 U10214 ( .B(n6751), .A(n6748), .S(n8520), .Y(n6755) );
  MUX2X1 U10215 ( .B(n6754), .A(n6739), .S(N17), .Y(n8299) );
  MUX2X1 U10216 ( .B(\RF[30][13] ), .A(\RF[31][13] ), .S(n8389), .Y(n6759) );
  MUX2X1 U10217 ( .B(\RF[28][13] ), .A(\RF[29][13] ), .S(n8389), .Y(n6758) );
  MUX2X1 U10218 ( .B(\RF[26][13] ), .A(\RF[27][13] ), .S(n8389), .Y(n6762) );
  MUX2X1 U10219 ( .B(\RF[24][13] ), .A(\RF[25][13] ), .S(n8389), .Y(n6761) );
  MUX2X1 U10220 ( .B(n6760), .A(n6757), .S(n8519), .Y(n6771) );
  MUX2X1 U10221 ( .B(\RF[22][13] ), .A(\RF[23][13] ), .S(n8389), .Y(n6765) );
  MUX2X1 U10222 ( .B(\RF[20][13] ), .A(\RF[21][13] ), .S(n8389), .Y(n6764) );
  MUX2X1 U10223 ( .B(\RF[18][13] ), .A(\RF[19][13] ), .S(n8389), .Y(n6768) );
  MUX2X1 U10224 ( .B(\RF[16][13] ), .A(\RF[17][13] ), .S(n8389), .Y(n6767) );
  MUX2X1 U10225 ( .B(n6766), .A(n6763), .S(n8520), .Y(n6770) );
  MUX2X1 U10226 ( .B(\RF[14][13] ), .A(\RF[15][13] ), .S(n8389), .Y(n6774) );
  MUX2X1 U10227 ( .B(\RF[12][13] ), .A(\RF[13][13] ), .S(n8389), .Y(n6773) );
  MUX2X1 U10228 ( .B(\RF[10][13] ), .A(\RF[11][13] ), .S(n8389), .Y(n6777) );
  MUX2X1 U10229 ( .B(\RF[8][13] ), .A(\RF[9][13] ), .S(n8389), .Y(n6776) );
  MUX2X1 U10230 ( .B(n6775), .A(n6772), .S(N15), .Y(n6786) );
  MUX2X1 U10231 ( .B(\RF[6][13] ), .A(\RF[7][13] ), .S(n8390), .Y(n6780) );
  MUX2X1 U10232 ( .B(\RF[4][13] ), .A(\RF[5][13] ), .S(n8390), .Y(n6779) );
  MUX2X1 U10233 ( .B(\RF[2][13] ), .A(\RF[3][13] ), .S(n8390), .Y(n6783) );
  MUX2X1 U10234 ( .B(\RF[0][13] ), .A(\RF[1][13] ), .S(n8390), .Y(n6782) );
  MUX2X1 U10235 ( .B(n6781), .A(n6778), .S(n8525), .Y(n6785) );
  MUX2X1 U10236 ( .B(n6784), .A(n6769), .S(N17), .Y(n8300) );
  MUX2X1 U10237 ( .B(\RF[30][14] ), .A(\RF[31][14] ), .S(n8390), .Y(n6789) );
  MUX2X1 U10238 ( .B(\RF[28][14] ), .A(\RF[29][14] ), .S(n8390), .Y(n6788) );
  MUX2X1 U10239 ( .B(\RF[26][14] ), .A(\RF[27][14] ), .S(n8390), .Y(n6792) );
  MUX2X1 U10240 ( .B(\RF[24][14] ), .A(\RF[25][14] ), .S(n8390), .Y(n6791) );
  MUX2X1 U10241 ( .B(n6790), .A(n6787), .S(n8530), .Y(n6801) );
  MUX2X1 U10242 ( .B(\RF[22][14] ), .A(\RF[23][14] ), .S(n8390), .Y(n6795) );
  MUX2X1 U10243 ( .B(\RF[20][14] ), .A(\RF[21][14] ), .S(n8390), .Y(n6794) );
  MUX2X1 U10244 ( .B(\RF[18][14] ), .A(\RF[19][14] ), .S(n8390), .Y(n6798) );
  MUX2X1 U10245 ( .B(\RF[16][14] ), .A(\RF[17][14] ), .S(n8390), .Y(n6797) );
  MUX2X1 U10246 ( .B(n6796), .A(n6793), .S(n8522), .Y(n6800) );
  MUX2X1 U10247 ( .B(\RF[14][14] ), .A(\RF[15][14] ), .S(n8391), .Y(n6804) );
  MUX2X1 U10248 ( .B(\RF[12][14] ), .A(\RF[13][14] ), .S(n8391), .Y(n6803) );
  MUX2X1 U10249 ( .B(\RF[10][14] ), .A(\RF[11][14] ), .S(n8391), .Y(n6807) );
  MUX2X1 U10250 ( .B(\RF[8][14] ), .A(\RF[9][14] ), .S(n8391), .Y(n6806) );
  MUX2X1 U10251 ( .B(n6805), .A(n6802), .S(n8531), .Y(n6816) );
  MUX2X1 U10252 ( .B(\RF[6][14] ), .A(\RF[7][14] ), .S(n8391), .Y(n6810) );
  MUX2X1 U10253 ( .B(\RF[4][14] ), .A(\RF[5][14] ), .S(n8391), .Y(n6809) );
  MUX2X1 U10254 ( .B(\RF[2][14] ), .A(\RF[3][14] ), .S(n8391), .Y(n6813) );
  MUX2X1 U10255 ( .B(\RF[0][14] ), .A(\RF[1][14] ), .S(n8391), .Y(n6812) );
  MUX2X1 U10256 ( .B(n6811), .A(n6808), .S(n8526), .Y(n6815) );
  MUX2X1 U10257 ( .B(n6814), .A(n6799), .S(N17), .Y(n8301) );
  MUX2X1 U10258 ( .B(\RF[30][15] ), .A(\RF[31][15] ), .S(n8391), .Y(n6819) );
  MUX2X1 U10259 ( .B(\RF[28][15] ), .A(\RF[29][15] ), .S(n8391), .Y(n6818) );
  MUX2X1 U10260 ( .B(\RF[26][15] ), .A(\RF[27][15] ), .S(n8391), .Y(n6822) );
  MUX2X1 U10261 ( .B(\RF[24][15] ), .A(\RF[25][15] ), .S(n8391), .Y(n6821) );
  MUX2X1 U10262 ( .B(n6820), .A(n6817), .S(n8528), .Y(n6831) );
  MUX2X1 U10263 ( .B(\RF[22][15] ), .A(\RF[23][15] ), .S(n8392), .Y(n6825) );
  MUX2X1 U10264 ( .B(\RF[20][15] ), .A(\RF[21][15] ), .S(n8392), .Y(n6824) );
  MUX2X1 U10265 ( .B(\RF[18][15] ), .A(\RF[19][15] ), .S(n8392), .Y(n6828) );
  MUX2X1 U10266 ( .B(\RF[16][15] ), .A(\RF[17][15] ), .S(n8392), .Y(n6827) );
  MUX2X1 U10267 ( .B(n6826), .A(n6823), .S(n8532), .Y(n6830) );
  MUX2X1 U10268 ( .B(\RF[14][15] ), .A(\RF[15][15] ), .S(n8392), .Y(n6834) );
  MUX2X1 U10269 ( .B(\RF[12][15] ), .A(\RF[13][15] ), .S(n8392), .Y(n6833) );
  MUX2X1 U10270 ( .B(\RF[10][15] ), .A(\RF[11][15] ), .S(n8392), .Y(n6837) );
  MUX2X1 U10271 ( .B(\RF[8][15] ), .A(\RF[9][15] ), .S(n8392), .Y(n6836) );
  MUX2X1 U10272 ( .B(n6835), .A(n6832), .S(n8533), .Y(n6846) );
  MUX2X1 U10273 ( .B(\RF[6][15] ), .A(\RF[7][15] ), .S(n8392), .Y(n6840) );
  MUX2X1 U10274 ( .B(\RF[4][15] ), .A(\RF[5][15] ), .S(n8392), .Y(n6839) );
  MUX2X1 U10275 ( .B(\RF[2][15] ), .A(\RF[3][15] ), .S(n8392), .Y(n6843) );
  MUX2X1 U10276 ( .B(\RF[0][15] ), .A(\RF[1][15] ), .S(n8392), .Y(n6842) );
  MUX2X1 U10277 ( .B(n6841), .A(n6838), .S(n8517), .Y(n6845) );
  MUX2X1 U10278 ( .B(n6844), .A(n6829), .S(N17), .Y(n8302) );
  MUX2X1 U10279 ( .B(\RF[30][16] ), .A(\RF[31][16] ), .S(n8393), .Y(n6849) );
  MUX2X1 U10280 ( .B(\RF[28][16] ), .A(\RF[29][16] ), .S(n8393), .Y(n6848) );
  MUX2X1 U10281 ( .B(\RF[26][16] ), .A(\RF[27][16] ), .S(n8393), .Y(n6852) );
  MUX2X1 U10282 ( .B(\RF[24][16] ), .A(\RF[25][16] ), .S(n8393), .Y(n6851) );
  MUX2X1 U10283 ( .B(n6850), .A(n6847), .S(n8521), .Y(n6861) );
  MUX2X1 U10284 ( .B(\RF[22][16] ), .A(\RF[23][16] ), .S(n8393), .Y(n6855) );
  MUX2X1 U10285 ( .B(\RF[20][16] ), .A(\RF[21][16] ), .S(n8393), .Y(n6854) );
  MUX2X1 U10286 ( .B(\RF[18][16] ), .A(\RF[19][16] ), .S(n8393), .Y(n6858) );
  MUX2X1 U10287 ( .B(\RF[16][16] ), .A(\RF[17][16] ), .S(n8393), .Y(n6857) );
  MUX2X1 U10288 ( .B(n6856), .A(n6853), .S(n8521), .Y(n6860) );
  MUX2X1 U10289 ( .B(\RF[14][16] ), .A(\RF[15][16] ), .S(n8393), .Y(n6864) );
  MUX2X1 U10290 ( .B(\RF[12][16] ), .A(\RF[13][16] ), .S(n8393), .Y(n6863) );
  MUX2X1 U10291 ( .B(\RF[10][16] ), .A(\RF[11][16] ), .S(n8393), .Y(n6867) );
  MUX2X1 U10292 ( .B(\RF[8][16] ), .A(\RF[9][16] ), .S(n8393), .Y(n6866) );
  MUX2X1 U10293 ( .B(n6865), .A(n6862), .S(n8521), .Y(n6876) );
  MUX2X1 U10294 ( .B(\RF[6][16] ), .A(\RF[7][16] ), .S(n8394), .Y(n6870) );
  MUX2X1 U10295 ( .B(\RF[4][16] ), .A(\RF[5][16] ), .S(n8394), .Y(n6869) );
  MUX2X1 U10296 ( .B(\RF[2][16] ), .A(\RF[3][16] ), .S(n8394), .Y(n6873) );
  MUX2X1 U10297 ( .B(\RF[0][16] ), .A(\RF[1][16] ), .S(n8394), .Y(n6872) );
  MUX2X1 U10298 ( .B(n6871), .A(n6868), .S(n8521), .Y(n6875) );
  MUX2X1 U10299 ( .B(n6874), .A(n6859), .S(N17), .Y(n8303) );
  MUX2X1 U10300 ( .B(\RF[30][17] ), .A(\RF[31][17] ), .S(n8394), .Y(n6879) );
  MUX2X1 U10301 ( .B(\RF[28][17] ), .A(\RF[29][17] ), .S(n8394), .Y(n6878) );
  MUX2X1 U10302 ( .B(\RF[26][17] ), .A(\RF[27][17] ), .S(n8394), .Y(n6882) );
  MUX2X1 U10303 ( .B(\RF[24][17] ), .A(\RF[25][17] ), .S(n8394), .Y(n6881) );
  MUX2X1 U10304 ( .B(n6880), .A(n6877), .S(n8521), .Y(n6891) );
  MUX2X1 U10305 ( .B(\RF[22][17] ), .A(\RF[23][17] ), .S(n8394), .Y(n6885) );
  MUX2X1 U10306 ( .B(\RF[20][17] ), .A(\RF[21][17] ), .S(n8394), .Y(n6884) );
  MUX2X1 U10307 ( .B(\RF[18][17] ), .A(\RF[19][17] ), .S(n8394), .Y(n6888) );
  MUX2X1 U10308 ( .B(\RF[16][17] ), .A(\RF[17][17] ), .S(n8394), .Y(n6887) );
  MUX2X1 U10309 ( .B(n6886), .A(n6883), .S(n8521), .Y(n6890) );
  MUX2X1 U10310 ( .B(\RF[14][17] ), .A(\RF[15][17] ), .S(n8395), .Y(n6894) );
  MUX2X1 U10311 ( .B(\RF[12][17] ), .A(\RF[13][17] ), .S(n8395), .Y(n6893) );
  MUX2X1 U10312 ( .B(\RF[10][17] ), .A(\RF[11][17] ), .S(n8395), .Y(n6897) );
  MUX2X1 U10313 ( .B(\RF[8][17] ), .A(\RF[9][17] ), .S(n8395), .Y(n6896) );
  MUX2X1 U10314 ( .B(n6895), .A(n6892), .S(n8521), .Y(n6906) );
  MUX2X1 U10315 ( .B(\RF[6][17] ), .A(\RF[7][17] ), .S(n8395), .Y(n6900) );
  MUX2X1 U10316 ( .B(\RF[4][17] ), .A(\RF[5][17] ), .S(n8395), .Y(n6899) );
  MUX2X1 U10317 ( .B(\RF[2][17] ), .A(\RF[3][17] ), .S(n8395), .Y(n6903) );
  MUX2X1 U10318 ( .B(\RF[0][17] ), .A(\RF[1][17] ), .S(n8395), .Y(n6902) );
  MUX2X1 U10319 ( .B(n6901), .A(n6898), .S(n8521), .Y(n6905) );
  MUX2X1 U10320 ( .B(n6904), .A(n6889), .S(N17), .Y(n8304) );
  MUX2X1 U10321 ( .B(\RF[30][18] ), .A(\RF[31][18] ), .S(n8395), .Y(n6909) );
  MUX2X1 U10322 ( .B(\RF[28][18] ), .A(\RF[29][18] ), .S(n8395), .Y(n6908) );
  MUX2X1 U10323 ( .B(\RF[26][18] ), .A(\RF[27][18] ), .S(n8395), .Y(n6912) );
  MUX2X1 U10324 ( .B(\RF[24][18] ), .A(\RF[25][18] ), .S(n8395), .Y(n6911) );
  MUX2X1 U10325 ( .B(n6910), .A(n6907), .S(n8521), .Y(n6921) );
  MUX2X1 U10326 ( .B(\RF[22][18] ), .A(\RF[23][18] ), .S(n8396), .Y(n6915) );
  MUX2X1 U10327 ( .B(\RF[20][18] ), .A(\RF[21][18] ), .S(n8396), .Y(n6914) );
  MUX2X1 U10328 ( .B(\RF[18][18] ), .A(\RF[19][18] ), .S(n8396), .Y(n6918) );
  MUX2X1 U10329 ( .B(\RF[16][18] ), .A(\RF[17][18] ), .S(n8396), .Y(n6917) );
  MUX2X1 U10330 ( .B(n6916), .A(n6913), .S(n8521), .Y(n6920) );
  MUX2X1 U10331 ( .B(\RF[14][18] ), .A(\RF[15][18] ), .S(n8396), .Y(n6924) );
  MUX2X1 U10332 ( .B(\RF[12][18] ), .A(\RF[13][18] ), .S(n8396), .Y(n6923) );
  MUX2X1 U10333 ( .B(\RF[10][18] ), .A(\RF[11][18] ), .S(n8396), .Y(n6927) );
  MUX2X1 U10334 ( .B(\RF[8][18] ), .A(\RF[9][18] ), .S(n8396), .Y(n6926) );
  MUX2X1 U10335 ( .B(n6925), .A(n6922), .S(n8521), .Y(n6936) );
  MUX2X1 U10336 ( .B(\RF[6][18] ), .A(\RF[7][18] ), .S(n8396), .Y(n6930) );
  MUX2X1 U10337 ( .B(\RF[4][18] ), .A(\RF[5][18] ), .S(n8396), .Y(n6929) );
  MUX2X1 U10338 ( .B(\RF[2][18] ), .A(\RF[3][18] ), .S(n8396), .Y(n6933) );
  MUX2X1 U10339 ( .B(\RF[0][18] ), .A(\RF[1][18] ), .S(n8396), .Y(n6932) );
  MUX2X1 U10340 ( .B(n6931), .A(n6928), .S(n8521), .Y(n6935) );
  MUX2X1 U10341 ( .B(n6934), .A(n6919), .S(N17), .Y(n8305) );
  MUX2X1 U10342 ( .B(\RF[30][19] ), .A(\RF[31][19] ), .S(n8397), .Y(n6939) );
  MUX2X1 U10343 ( .B(\RF[28][19] ), .A(\RF[29][19] ), .S(n8397), .Y(n6938) );
  MUX2X1 U10344 ( .B(\RF[26][19] ), .A(\RF[27][19] ), .S(n8397), .Y(n6942) );
  MUX2X1 U10345 ( .B(\RF[24][19] ), .A(\RF[25][19] ), .S(n8397), .Y(n6941) );
  MUX2X1 U10346 ( .B(n6940), .A(n6937), .S(n8522), .Y(n6951) );
  MUX2X1 U10347 ( .B(\RF[22][19] ), .A(\RF[23][19] ), .S(n8397), .Y(n6945) );
  MUX2X1 U10348 ( .B(\RF[20][19] ), .A(\RF[21][19] ), .S(n8397), .Y(n6944) );
  MUX2X1 U10349 ( .B(\RF[18][19] ), .A(\RF[19][19] ), .S(n8397), .Y(n6948) );
  MUX2X1 U10350 ( .B(\RF[16][19] ), .A(\RF[17][19] ), .S(n8397), .Y(n6947) );
  MUX2X1 U10351 ( .B(n6946), .A(n6943), .S(n8522), .Y(n6950) );
  MUX2X1 U10352 ( .B(\RF[14][19] ), .A(\RF[15][19] ), .S(n8397), .Y(n6954) );
  MUX2X1 U10353 ( .B(\RF[12][19] ), .A(\RF[13][19] ), .S(n8397), .Y(n6953) );
  MUX2X1 U10354 ( .B(\RF[10][19] ), .A(\RF[11][19] ), .S(n8397), .Y(n6957) );
  MUX2X1 U10355 ( .B(\RF[8][19] ), .A(\RF[9][19] ), .S(n8397), .Y(n6956) );
  MUX2X1 U10356 ( .B(n6955), .A(n6952), .S(n8522), .Y(n6966) );
  MUX2X1 U10357 ( .B(\RF[6][19] ), .A(\RF[7][19] ), .S(n8398), .Y(n6960) );
  MUX2X1 U10358 ( .B(\RF[4][19] ), .A(\RF[5][19] ), .S(n8398), .Y(n6959) );
  MUX2X1 U10359 ( .B(\RF[2][19] ), .A(\RF[3][19] ), .S(n8398), .Y(n6963) );
  MUX2X1 U10360 ( .B(\RF[0][19] ), .A(\RF[1][19] ), .S(n8398), .Y(n6962) );
  MUX2X1 U10361 ( .B(n6961), .A(n6958), .S(n8522), .Y(n6965) );
  MUX2X1 U10362 ( .B(n6964), .A(n6949), .S(N17), .Y(n8306) );
  MUX2X1 U10363 ( .B(\RF[30][20] ), .A(\RF[31][20] ), .S(n8398), .Y(n6969) );
  MUX2X1 U10364 ( .B(\RF[28][20] ), .A(\RF[29][20] ), .S(n8398), .Y(n6968) );
  MUX2X1 U10365 ( .B(\RF[26][20] ), .A(\RF[27][20] ), .S(n8398), .Y(n6972) );
  MUX2X1 U10366 ( .B(\RF[24][20] ), .A(\RF[25][20] ), .S(n8398), .Y(n6971) );
  MUX2X1 U10367 ( .B(n6970), .A(n6967), .S(n8522), .Y(n6981) );
  MUX2X1 U10368 ( .B(\RF[22][20] ), .A(\RF[23][20] ), .S(n8398), .Y(n6975) );
  MUX2X1 U10369 ( .B(\RF[20][20] ), .A(\RF[21][20] ), .S(n8398), .Y(n6974) );
  MUX2X1 U10370 ( .B(\RF[18][20] ), .A(\RF[19][20] ), .S(n8398), .Y(n6978) );
  MUX2X1 U10371 ( .B(\RF[16][20] ), .A(\RF[17][20] ), .S(n8398), .Y(n6977) );
  MUX2X1 U10372 ( .B(n6976), .A(n6973), .S(n8522), .Y(n6980) );
  MUX2X1 U10373 ( .B(\RF[14][20] ), .A(\RF[15][20] ), .S(n8399), .Y(n6984) );
  MUX2X1 U10374 ( .B(\RF[12][20] ), .A(\RF[13][20] ), .S(n8399), .Y(n6983) );
  MUX2X1 U10375 ( .B(\RF[10][20] ), .A(\RF[11][20] ), .S(n8399), .Y(n6987) );
  MUX2X1 U10376 ( .B(\RF[8][20] ), .A(\RF[9][20] ), .S(n8399), .Y(n6986) );
  MUX2X1 U10377 ( .B(n6985), .A(n6982), .S(n8522), .Y(n6996) );
  MUX2X1 U10378 ( .B(\RF[6][20] ), .A(\RF[7][20] ), .S(n8399), .Y(n6990) );
  MUX2X1 U10379 ( .B(\RF[4][20] ), .A(\RF[5][20] ), .S(n8399), .Y(n6989) );
  MUX2X1 U10380 ( .B(\RF[2][20] ), .A(\RF[3][20] ), .S(n8399), .Y(n6993) );
  MUX2X1 U10381 ( .B(\RF[0][20] ), .A(\RF[1][20] ), .S(n8399), .Y(n6992) );
  MUX2X1 U10382 ( .B(n6991), .A(n6988), .S(n8522), .Y(n6995) );
  MUX2X1 U10383 ( .B(n6994), .A(n6979), .S(N17), .Y(n8307) );
  MUX2X1 U10384 ( .B(\RF[30][21] ), .A(\RF[31][21] ), .S(n8399), .Y(n6999) );
  MUX2X1 U10385 ( .B(\RF[28][21] ), .A(\RF[29][21] ), .S(n8399), .Y(n6998) );
  MUX2X1 U10386 ( .B(\RF[26][21] ), .A(\RF[27][21] ), .S(n8399), .Y(n7002) );
  MUX2X1 U10387 ( .B(\RF[24][21] ), .A(\RF[25][21] ), .S(n8399), .Y(n7001) );
  MUX2X1 U10388 ( .B(n7000), .A(n6997), .S(n8522), .Y(n7011) );
  MUX2X1 U10389 ( .B(\RF[22][21] ), .A(\RF[23][21] ), .S(n8400), .Y(n7005) );
  MUX2X1 U10390 ( .B(\RF[20][21] ), .A(\RF[21][21] ), .S(n8400), .Y(n7004) );
  MUX2X1 U10391 ( .B(\RF[18][21] ), .A(\RF[19][21] ), .S(n8400), .Y(n7008) );
  MUX2X1 U10392 ( .B(\RF[16][21] ), .A(\RF[17][21] ), .S(n8400), .Y(n7007) );
  MUX2X1 U10393 ( .B(n7006), .A(n7003), .S(n8522), .Y(n7010) );
  MUX2X1 U10394 ( .B(\RF[14][21] ), .A(\RF[15][21] ), .S(n8400), .Y(n7014) );
  MUX2X1 U10395 ( .B(\RF[12][21] ), .A(\RF[13][21] ), .S(n8400), .Y(n7013) );
  MUX2X1 U10396 ( .B(\RF[10][21] ), .A(\RF[11][21] ), .S(n8400), .Y(n7017) );
  MUX2X1 U10397 ( .B(\RF[8][21] ), .A(\RF[9][21] ), .S(n8400), .Y(n7016) );
  MUX2X1 U10398 ( .B(n7015), .A(n7012), .S(n8522), .Y(n7026) );
  MUX2X1 U10399 ( .B(\RF[6][21] ), .A(\RF[7][21] ), .S(n8400), .Y(n7020) );
  MUX2X1 U10400 ( .B(\RF[4][21] ), .A(\RF[5][21] ), .S(n8400), .Y(n7019) );
  MUX2X1 U10401 ( .B(\RF[2][21] ), .A(\RF[3][21] ), .S(n8400), .Y(n7023) );
  MUX2X1 U10402 ( .B(\RF[0][21] ), .A(\RF[1][21] ), .S(n8400), .Y(n7022) );
  MUX2X1 U10403 ( .B(n7021), .A(n7018), .S(n8522), .Y(n7025) );
  MUX2X1 U10404 ( .B(n7024), .A(n7009), .S(N17), .Y(n8308) );
  MUX2X1 U10405 ( .B(\RF[30][22] ), .A(\RF[31][22] ), .S(n8401), .Y(n7029) );
  MUX2X1 U10406 ( .B(\RF[28][22] ), .A(\RF[29][22] ), .S(n8401), .Y(n7028) );
  MUX2X1 U10407 ( .B(\RF[26][22] ), .A(\RF[27][22] ), .S(n8401), .Y(n7032) );
  MUX2X1 U10408 ( .B(\RF[24][22] ), .A(\RF[25][22] ), .S(n8401), .Y(n7031) );
  MUX2X1 U10409 ( .B(n7030), .A(n7027), .S(n8523), .Y(n7041) );
  MUX2X1 U10410 ( .B(\RF[22][22] ), .A(\RF[23][22] ), .S(n8401), .Y(n7035) );
  MUX2X1 U10411 ( .B(\RF[20][22] ), .A(\RF[21][22] ), .S(n8401), .Y(n7034) );
  MUX2X1 U10412 ( .B(\RF[18][22] ), .A(\RF[19][22] ), .S(n8401), .Y(n7038) );
  MUX2X1 U10413 ( .B(\RF[16][22] ), .A(\RF[17][22] ), .S(n8401), .Y(n7037) );
  MUX2X1 U10414 ( .B(n7036), .A(n7033), .S(n8523), .Y(n7040) );
  MUX2X1 U10415 ( .B(\RF[14][22] ), .A(\RF[15][22] ), .S(n8401), .Y(n7044) );
  MUX2X1 U10416 ( .B(\RF[12][22] ), .A(\RF[13][22] ), .S(n8401), .Y(n7043) );
  MUX2X1 U10417 ( .B(\RF[10][22] ), .A(\RF[11][22] ), .S(n8401), .Y(n7047) );
  MUX2X1 U10418 ( .B(\RF[8][22] ), .A(\RF[9][22] ), .S(n8401), .Y(n7046) );
  MUX2X1 U10419 ( .B(n7045), .A(n7042), .S(n8523), .Y(n7056) );
  MUX2X1 U10420 ( .B(\RF[6][22] ), .A(\RF[7][22] ), .S(n8402), .Y(n7050) );
  MUX2X1 U10421 ( .B(\RF[4][22] ), .A(\RF[5][22] ), .S(n8402), .Y(n7049) );
  MUX2X1 U10422 ( .B(\RF[2][22] ), .A(\RF[3][22] ), .S(n8402), .Y(n7053) );
  MUX2X1 U10423 ( .B(\RF[0][22] ), .A(\RF[1][22] ), .S(n8402), .Y(n7052) );
  MUX2X1 U10424 ( .B(n7051), .A(n7048), .S(n8523), .Y(n7055) );
  MUX2X1 U10425 ( .B(n7054), .A(n7039), .S(N17), .Y(n8309) );
  MUX2X1 U10426 ( .B(\RF[30][23] ), .A(\RF[31][23] ), .S(n8402), .Y(n7059) );
  MUX2X1 U10427 ( .B(\RF[28][23] ), .A(\RF[29][23] ), .S(n8402), .Y(n7058) );
  MUX2X1 U10428 ( .B(\RF[26][23] ), .A(\RF[27][23] ), .S(n8402), .Y(n7062) );
  MUX2X1 U10429 ( .B(\RF[24][23] ), .A(\RF[25][23] ), .S(n8402), .Y(n7061) );
  MUX2X1 U10430 ( .B(n7060), .A(n7057), .S(n8523), .Y(n7071) );
  MUX2X1 U10431 ( .B(\RF[22][23] ), .A(\RF[23][23] ), .S(n8402), .Y(n7065) );
  MUX2X1 U10432 ( .B(\RF[20][23] ), .A(\RF[21][23] ), .S(n8402), .Y(n7064) );
  MUX2X1 U10433 ( .B(\RF[18][23] ), .A(\RF[19][23] ), .S(n8402), .Y(n7068) );
  MUX2X1 U10434 ( .B(\RF[16][23] ), .A(\RF[17][23] ), .S(n8402), .Y(n7067) );
  MUX2X1 U10435 ( .B(n7066), .A(n7063), .S(n8523), .Y(n7070) );
  MUX2X1 U10436 ( .B(\RF[14][23] ), .A(\RF[15][23] ), .S(n8403), .Y(n7074) );
  MUX2X1 U10437 ( .B(\RF[12][23] ), .A(\RF[13][23] ), .S(n8403), .Y(n7073) );
  MUX2X1 U10438 ( .B(\RF[10][23] ), .A(\RF[11][23] ), .S(n8403), .Y(n7077) );
  MUX2X1 U10439 ( .B(\RF[8][23] ), .A(\RF[9][23] ), .S(n8403), .Y(n7076) );
  MUX2X1 U10440 ( .B(n7075), .A(n7072), .S(n8523), .Y(n7086) );
  MUX2X1 U10441 ( .B(\RF[6][23] ), .A(\RF[7][23] ), .S(n8403), .Y(n7080) );
  MUX2X1 U10442 ( .B(\RF[4][23] ), .A(\RF[5][23] ), .S(n8403), .Y(n7079) );
  MUX2X1 U10443 ( .B(\RF[2][23] ), .A(\RF[3][23] ), .S(n8403), .Y(n7083) );
  MUX2X1 U10444 ( .B(\RF[0][23] ), .A(\RF[1][23] ), .S(n8403), .Y(n7082) );
  MUX2X1 U10445 ( .B(n7081), .A(n7078), .S(n8523), .Y(n7085) );
  MUX2X1 U10446 ( .B(n7084), .A(n7069), .S(N17), .Y(n8310) );
  MUX2X1 U10447 ( .B(\RF[30][24] ), .A(\RF[31][24] ), .S(n8403), .Y(n7089) );
  MUX2X1 U10448 ( .B(\RF[28][24] ), .A(\RF[29][24] ), .S(n8403), .Y(n7088) );
  MUX2X1 U10449 ( .B(\RF[26][24] ), .A(\RF[27][24] ), .S(n8403), .Y(n7092) );
  MUX2X1 U10450 ( .B(\RF[24][24] ), .A(\RF[25][24] ), .S(n8403), .Y(n7091) );
  MUX2X1 U10451 ( .B(n7090), .A(n7087), .S(n8523), .Y(n7101) );
  MUX2X1 U10452 ( .B(\RF[22][24] ), .A(\RF[23][24] ), .S(n8404), .Y(n7095) );
  MUX2X1 U10453 ( .B(\RF[20][24] ), .A(\RF[21][24] ), .S(n8404), .Y(n7094) );
  MUX2X1 U10454 ( .B(\RF[18][24] ), .A(\RF[19][24] ), .S(n8404), .Y(n7098) );
  MUX2X1 U10455 ( .B(\RF[16][24] ), .A(\RF[17][24] ), .S(n8404), .Y(n7097) );
  MUX2X1 U10456 ( .B(n7096), .A(n7093), .S(n8523), .Y(n7100) );
  MUX2X1 U10457 ( .B(\RF[14][24] ), .A(\RF[15][24] ), .S(n8404), .Y(n7104) );
  MUX2X1 U10458 ( .B(\RF[12][24] ), .A(\RF[13][24] ), .S(n8404), .Y(n7103) );
  MUX2X1 U10459 ( .B(\RF[10][24] ), .A(\RF[11][24] ), .S(n8404), .Y(n7107) );
  MUX2X1 U10460 ( .B(\RF[8][24] ), .A(\RF[9][24] ), .S(n8404), .Y(n7106) );
  MUX2X1 U10461 ( .B(n7105), .A(n7102), .S(n8523), .Y(n7116) );
  MUX2X1 U10462 ( .B(\RF[6][24] ), .A(\RF[7][24] ), .S(n8404), .Y(n7110) );
  MUX2X1 U10463 ( .B(\RF[4][24] ), .A(\RF[5][24] ), .S(n8404), .Y(n7109) );
  MUX2X1 U10464 ( .B(\RF[2][24] ), .A(\RF[3][24] ), .S(n8404), .Y(n7113) );
  MUX2X1 U10465 ( .B(\RF[0][24] ), .A(\RF[1][24] ), .S(n8404), .Y(n7112) );
  MUX2X1 U10466 ( .B(n7111), .A(n7108), .S(n8523), .Y(n7115) );
  MUX2X1 U10467 ( .B(n7114), .A(n7099), .S(N17), .Y(n8311) );
  MUX2X1 U10468 ( .B(\RF[30][25] ), .A(\RF[31][25] ), .S(n8405), .Y(n7119) );
  MUX2X1 U10469 ( .B(\RF[28][25] ), .A(\RF[29][25] ), .S(n8405), .Y(n7118) );
  MUX2X1 U10470 ( .B(\RF[26][25] ), .A(\RF[27][25] ), .S(n8405), .Y(n7122) );
  MUX2X1 U10471 ( .B(\RF[24][25] ), .A(\RF[25][25] ), .S(n8405), .Y(n7121) );
  MUX2X1 U10472 ( .B(n7120), .A(n7117), .S(n8524), .Y(n7131) );
  MUX2X1 U10473 ( .B(\RF[22][25] ), .A(\RF[23][25] ), .S(n8405), .Y(n7125) );
  MUX2X1 U10474 ( .B(\RF[20][25] ), .A(\RF[21][25] ), .S(n8405), .Y(n7124) );
  MUX2X1 U10475 ( .B(\RF[18][25] ), .A(\RF[19][25] ), .S(n8405), .Y(n7128) );
  MUX2X1 U10476 ( .B(\RF[16][25] ), .A(\RF[17][25] ), .S(n8405), .Y(n7127) );
  MUX2X1 U10477 ( .B(n7126), .A(n7123), .S(n8524), .Y(n7130) );
  MUX2X1 U10478 ( .B(\RF[14][25] ), .A(\RF[15][25] ), .S(n8405), .Y(n7134) );
  MUX2X1 U10479 ( .B(\RF[12][25] ), .A(\RF[13][25] ), .S(n8405), .Y(n7133) );
  MUX2X1 U10480 ( .B(\RF[10][25] ), .A(\RF[11][25] ), .S(n8405), .Y(n7137) );
  MUX2X1 U10481 ( .B(\RF[8][25] ), .A(\RF[9][25] ), .S(n8405), .Y(n7136) );
  MUX2X1 U10482 ( .B(n7135), .A(n7132), .S(n8524), .Y(n7146) );
  MUX2X1 U10483 ( .B(\RF[6][25] ), .A(\RF[7][25] ), .S(n8406), .Y(n7140) );
  MUX2X1 U10484 ( .B(\RF[4][25] ), .A(\RF[5][25] ), .S(n8406), .Y(n7139) );
  MUX2X1 U10485 ( .B(\RF[2][25] ), .A(\RF[3][25] ), .S(n8406), .Y(n7143) );
  MUX2X1 U10486 ( .B(\RF[0][25] ), .A(\RF[1][25] ), .S(n8406), .Y(n7142) );
  MUX2X1 U10487 ( .B(n7141), .A(n7138), .S(n8524), .Y(n7145) );
  MUX2X1 U10488 ( .B(n7144), .A(n7129), .S(N17), .Y(n8312) );
  MUX2X1 U10489 ( .B(\RF[30][26] ), .A(\RF[31][26] ), .S(n8406), .Y(n7149) );
  MUX2X1 U10490 ( .B(\RF[28][26] ), .A(\RF[29][26] ), .S(n8406), .Y(n7148) );
  MUX2X1 U10491 ( .B(\RF[26][26] ), .A(\RF[27][26] ), .S(n8406), .Y(n7152) );
  MUX2X1 U10492 ( .B(\RF[24][26] ), .A(\RF[25][26] ), .S(n8406), .Y(n7151) );
  MUX2X1 U10493 ( .B(n7150), .A(n7147), .S(n8524), .Y(n7161) );
  MUX2X1 U10494 ( .B(\RF[22][26] ), .A(\RF[23][26] ), .S(n8406), .Y(n7155) );
  MUX2X1 U10495 ( .B(\RF[20][26] ), .A(\RF[21][26] ), .S(n8406), .Y(n7154) );
  MUX2X1 U10496 ( .B(\RF[18][26] ), .A(\RF[19][26] ), .S(n8406), .Y(n7158) );
  MUX2X1 U10497 ( .B(\RF[16][26] ), .A(\RF[17][26] ), .S(n8406), .Y(n7157) );
  MUX2X1 U10498 ( .B(n7156), .A(n7153), .S(n8524), .Y(n7160) );
  MUX2X1 U10499 ( .B(\RF[14][26] ), .A(\RF[15][26] ), .S(n8407), .Y(n7164) );
  MUX2X1 U10500 ( .B(\RF[12][26] ), .A(\RF[13][26] ), .S(n8407), .Y(n7163) );
  MUX2X1 U10501 ( .B(\RF[10][26] ), .A(\RF[11][26] ), .S(n8407), .Y(n7167) );
  MUX2X1 U10502 ( .B(\RF[8][26] ), .A(\RF[9][26] ), .S(n8407), .Y(n7166) );
  MUX2X1 U10503 ( .B(n7165), .A(n7162), .S(n8524), .Y(n7176) );
  MUX2X1 U10504 ( .B(\RF[6][26] ), .A(\RF[7][26] ), .S(n8407), .Y(n7170) );
  MUX2X1 U10505 ( .B(\RF[4][26] ), .A(\RF[5][26] ), .S(n8407), .Y(n7169) );
  MUX2X1 U10506 ( .B(\RF[2][26] ), .A(\RF[3][26] ), .S(n8407), .Y(n7173) );
  MUX2X1 U10507 ( .B(\RF[0][26] ), .A(\RF[1][26] ), .S(n8407), .Y(n7172) );
  MUX2X1 U10508 ( .B(n7171), .A(n7168), .S(n8524), .Y(n7175) );
  MUX2X1 U10509 ( .B(n7174), .A(n7159), .S(N17), .Y(n8313) );
  MUX2X1 U10510 ( .B(\RF[30][27] ), .A(\RF[31][27] ), .S(n8407), .Y(n7179) );
  MUX2X1 U10511 ( .B(\RF[28][27] ), .A(\RF[29][27] ), .S(n8407), .Y(n7178) );
  MUX2X1 U10512 ( .B(\RF[26][27] ), .A(\RF[27][27] ), .S(n8407), .Y(n7182) );
  MUX2X1 U10513 ( .B(\RF[24][27] ), .A(\RF[25][27] ), .S(n8407), .Y(n7181) );
  MUX2X1 U10514 ( .B(n7180), .A(n7177), .S(n8524), .Y(n7191) );
  MUX2X1 U10515 ( .B(\RF[22][27] ), .A(\RF[23][27] ), .S(n8408), .Y(n7185) );
  MUX2X1 U10516 ( .B(\RF[20][27] ), .A(\RF[21][27] ), .S(n8408), .Y(n7184) );
  MUX2X1 U10517 ( .B(\RF[18][27] ), .A(\RF[19][27] ), .S(n8408), .Y(n7188) );
  MUX2X1 U10518 ( .B(\RF[16][27] ), .A(\RF[17][27] ), .S(n8408), .Y(n7187) );
  MUX2X1 U10519 ( .B(n7186), .A(n7183), .S(n8524), .Y(n7190) );
  MUX2X1 U10520 ( .B(\RF[14][27] ), .A(\RF[15][27] ), .S(n8408), .Y(n7194) );
  MUX2X1 U10521 ( .B(\RF[12][27] ), .A(\RF[13][27] ), .S(n8408), .Y(n7193) );
  MUX2X1 U10522 ( .B(\RF[10][27] ), .A(\RF[11][27] ), .S(n8408), .Y(n7197) );
  MUX2X1 U10523 ( .B(\RF[8][27] ), .A(\RF[9][27] ), .S(n8408), .Y(n7196) );
  MUX2X1 U10524 ( .B(n7195), .A(n7192), .S(n8524), .Y(n7206) );
  MUX2X1 U10525 ( .B(\RF[6][27] ), .A(\RF[7][27] ), .S(n8408), .Y(n7200) );
  MUX2X1 U10526 ( .B(\RF[4][27] ), .A(\RF[5][27] ), .S(n8408), .Y(n7199) );
  MUX2X1 U10527 ( .B(\RF[2][27] ), .A(\RF[3][27] ), .S(n8408), .Y(n7203) );
  MUX2X1 U10528 ( .B(\RF[0][27] ), .A(\RF[1][27] ), .S(n8408), .Y(n7202) );
  MUX2X1 U10529 ( .B(n7201), .A(n7198), .S(n8524), .Y(n7205) );
  MUX2X1 U10530 ( .B(n7204), .A(n7189), .S(N17), .Y(n8314) );
  MUX2X1 U10531 ( .B(\RF[30][28] ), .A(\RF[31][28] ), .S(n8409), .Y(n7209) );
  MUX2X1 U10532 ( .B(\RF[28][28] ), .A(\RF[29][28] ), .S(n8409), .Y(n7208) );
  MUX2X1 U10533 ( .B(\RF[26][28] ), .A(\RF[27][28] ), .S(n8409), .Y(n7212) );
  MUX2X1 U10534 ( .B(\RF[24][28] ), .A(\RF[25][28] ), .S(n8409), .Y(n7211) );
  MUX2X1 U10535 ( .B(n7210), .A(n7207), .S(n8525), .Y(n7221) );
  MUX2X1 U10536 ( .B(\RF[22][28] ), .A(\RF[23][28] ), .S(n8409), .Y(n7215) );
  MUX2X1 U10537 ( .B(\RF[20][28] ), .A(\RF[21][28] ), .S(n8409), .Y(n7214) );
  MUX2X1 U10538 ( .B(\RF[18][28] ), .A(\RF[19][28] ), .S(n8409), .Y(n7218) );
  MUX2X1 U10539 ( .B(\RF[16][28] ), .A(\RF[17][28] ), .S(n8409), .Y(n7217) );
  MUX2X1 U10540 ( .B(n7216), .A(n7213), .S(n8525), .Y(n7220) );
  MUX2X1 U10541 ( .B(\RF[14][28] ), .A(\RF[15][28] ), .S(n8409), .Y(n7224) );
  MUX2X1 U10542 ( .B(\RF[12][28] ), .A(\RF[13][28] ), .S(n8409), .Y(n7223) );
  MUX2X1 U10543 ( .B(\RF[10][28] ), .A(\RF[11][28] ), .S(n8409), .Y(n7227) );
  MUX2X1 U10544 ( .B(\RF[8][28] ), .A(\RF[9][28] ), .S(n8409), .Y(n7226) );
  MUX2X1 U10545 ( .B(n7225), .A(n7222), .S(n8525), .Y(n7236) );
  MUX2X1 U10546 ( .B(\RF[6][28] ), .A(\RF[7][28] ), .S(n8410), .Y(n7230) );
  MUX2X1 U10547 ( .B(\RF[4][28] ), .A(\RF[5][28] ), .S(n8410), .Y(n7229) );
  MUX2X1 U10548 ( .B(\RF[2][28] ), .A(\RF[3][28] ), .S(n8410), .Y(n7233) );
  MUX2X1 U10549 ( .B(\RF[0][28] ), .A(\RF[1][28] ), .S(n8410), .Y(n7232) );
  MUX2X1 U10550 ( .B(n7231), .A(n7228), .S(n8525), .Y(n7235) );
  MUX2X1 U10551 ( .B(n7234), .A(n7219), .S(N17), .Y(n8315) );
  MUX2X1 U10552 ( .B(\RF[30][29] ), .A(\RF[31][29] ), .S(n8410), .Y(n7239) );
  MUX2X1 U10553 ( .B(\RF[28][29] ), .A(\RF[29][29] ), .S(n8410), .Y(n7238) );
  MUX2X1 U10554 ( .B(\RF[26][29] ), .A(\RF[27][29] ), .S(n8410), .Y(n7242) );
  MUX2X1 U10555 ( .B(\RF[24][29] ), .A(\RF[25][29] ), .S(n8410), .Y(n7241) );
  MUX2X1 U10556 ( .B(n7240), .A(n7237), .S(n8525), .Y(n7251) );
  MUX2X1 U10557 ( .B(\RF[22][29] ), .A(\RF[23][29] ), .S(n8410), .Y(n7245) );
  MUX2X1 U10558 ( .B(\RF[20][29] ), .A(\RF[21][29] ), .S(n8410), .Y(n7244) );
  MUX2X1 U10559 ( .B(\RF[18][29] ), .A(\RF[19][29] ), .S(n8410), .Y(n7248) );
  MUX2X1 U10560 ( .B(\RF[16][29] ), .A(\RF[17][29] ), .S(n8410), .Y(n7247) );
  MUX2X1 U10561 ( .B(n7246), .A(n7243), .S(n8525), .Y(n7250) );
  MUX2X1 U10562 ( .B(\RF[14][29] ), .A(\RF[15][29] ), .S(n8411), .Y(n7254) );
  MUX2X1 U10563 ( .B(\RF[12][29] ), .A(\RF[13][29] ), .S(n8411), .Y(n7253) );
  MUX2X1 U10564 ( .B(\RF[10][29] ), .A(\RF[11][29] ), .S(n8411), .Y(n7257) );
  MUX2X1 U10565 ( .B(\RF[8][29] ), .A(\RF[9][29] ), .S(n8411), .Y(n7256) );
  MUX2X1 U10566 ( .B(n7255), .A(n7252), .S(n8525), .Y(n7266) );
  MUX2X1 U10567 ( .B(\RF[6][29] ), .A(\RF[7][29] ), .S(n8411), .Y(n7260) );
  MUX2X1 U10568 ( .B(\RF[4][29] ), .A(\RF[5][29] ), .S(n8411), .Y(n7259) );
  MUX2X1 U10569 ( .B(\RF[2][29] ), .A(\RF[3][29] ), .S(n8411), .Y(n7263) );
  MUX2X1 U10570 ( .B(\RF[0][29] ), .A(\RF[1][29] ), .S(n8411), .Y(n7262) );
  MUX2X1 U10571 ( .B(n7261), .A(n7258), .S(n8525), .Y(n7265) );
  MUX2X1 U10572 ( .B(n7264), .A(n7249), .S(N17), .Y(n8316) );
  MUX2X1 U10573 ( .B(\RF[30][30] ), .A(\RF[31][30] ), .S(n8411), .Y(n7269) );
  MUX2X1 U10574 ( .B(\RF[28][30] ), .A(\RF[29][30] ), .S(n8411), .Y(n7268) );
  MUX2X1 U10575 ( .B(\RF[26][30] ), .A(\RF[27][30] ), .S(n8411), .Y(n7272) );
  MUX2X1 U10576 ( .B(\RF[24][30] ), .A(\RF[25][30] ), .S(n8411), .Y(n7271) );
  MUX2X1 U10577 ( .B(n7270), .A(n7267), .S(n8525), .Y(n7281) );
  MUX2X1 U10578 ( .B(\RF[22][30] ), .A(\RF[23][30] ), .S(n8412), .Y(n7275) );
  MUX2X1 U10579 ( .B(\RF[20][30] ), .A(\RF[21][30] ), .S(n8412), .Y(n7274) );
  MUX2X1 U10580 ( .B(\RF[18][30] ), .A(\RF[19][30] ), .S(n8412), .Y(n7278) );
  MUX2X1 U10581 ( .B(\RF[16][30] ), .A(\RF[17][30] ), .S(n8412), .Y(n7277) );
  MUX2X1 U10582 ( .B(n7276), .A(n7273), .S(n8525), .Y(n7280) );
  MUX2X1 U10583 ( .B(\RF[14][30] ), .A(\RF[15][30] ), .S(n8412), .Y(n7284) );
  MUX2X1 U10584 ( .B(\RF[12][30] ), .A(\RF[13][30] ), .S(n8412), .Y(n7283) );
  MUX2X1 U10585 ( .B(\RF[10][30] ), .A(\RF[11][30] ), .S(n8412), .Y(n7287) );
  MUX2X1 U10586 ( .B(\RF[8][30] ), .A(\RF[9][30] ), .S(n8412), .Y(n7286) );
  MUX2X1 U10587 ( .B(n7285), .A(n7282), .S(n8525), .Y(n7296) );
  MUX2X1 U10588 ( .B(\RF[6][30] ), .A(\RF[7][30] ), .S(n8412), .Y(n7290) );
  MUX2X1 U10589 ( .B(\RF[4][30] ), .A(\RF[5][30] ), .S(n8412), .Y(n7289) );
  MUX2X1 U10590 ( .B(\RF[2][30] ), .A(\RF[3][30] ), .S(n8412), .Y(n7293) );
  MUX2X1 U10591 ( .B(\RF[0][30] ), .A(\RF[1][30] ), .S(n8412), .Y(n7292) );
  MUX2X1 U10592 ( .B(n7291), .A(n7288), .S(n8525), .Y(n7295) );
  MUX2X1 U10593 ( .B(n7294), .A(n7279), .S(N17), .Y(n8317) );
  MUX2X1 U10594 ( .B(\RF[30][31] ), .A(\RF[31][31] ), .S(n8413), .Y(n7299) );
  MUX2X1 U10595 ( .B(\RF[28][31] ), .A(\RF[29][31] ), .S(n8413), .Y(n7298) );
  MUX2X1 U10596 ( .B(\RF[26][31] ), .A(\RF[27][31] ), .S(n8413), .Y(n7302) );
  MUX2X1 U10597 ( .B(\RF[24][31] ), .A(\RF[25][31] ), .S(n8413), .Y(n7301) );
  MUX2X1 U10598 ( .B(n7300), .A(n7297), .S(n8526), .Y(n7311) );
  MUX2X1 U10599 ( .B(\RF[22][31] ), .A(\RF[23][31] ), .S(n8413), .Y(n7305) );
  MUX2X1 U10600 ( .B(\RF[20][31] ), .A(\RF[21][31] ), .S(n8413), .Y(n7304) );
  MUX2X1 U10601 ( .B(\RF[18][31] ), .A(\RF[19][31] ), .S(n8413), .Y(n7308) );
  MUX2X1 U10602 ( .B(\RF[16][31] ), .A(\RF[17][31] ), .S(n8413), .Y(n7307) );
  MUX2X1 U10603 ( .B(n7306), .A(n7303), .S(n8526), .Y(n7310) );
  MUX2X1 U10604 ( .B(\RF[14][31] ), .A(\RF[15][31] ), .S(n8413), .Y(n7314) );
  MUX2X1 U10605 ( .B(\RF[12][31] ), .A(\RF[13][31] ), .S(n8413), .Y(n7313) );
  MUX2X1 U10606 ( .B(\RF[10][31] ), .A(\RF[11][31] ), .S(n8413), .Y(n7317) );
  MUX2X1 U10607 ( .B(\RF[8][31] ), .A(\RF[9][31] ), .S(n8413), .Y(n7316) );
  MUX2X1 U10608 ( .B(n7315), .A(n7312), .S(n8526), .Y(n7326) );
  MUX2X1 U10609 ( .B(\RF[6][31] ), .A(\RF[7][31] ), .S(n8414), .Y(n7320) );
  MUX2X1 U10610 ( .B(\RF[4][31] ), .A(\RF[5][31] ), .S(n8414), .Y(n7319) );
  MUX2X1 U10611 ( .B(\RF[2][31] ), .A(\RF[3][31] ), .S(n8414), .Y(n7323) );
  MUX2X1 U10612 ( .B(\RF[0][31] ), .A(\RF[1][31] ), .S(n8414), .Y(n7322) );
  MUX2X1 U10613 ( .B(n7321), .A(n7318), .S(n8526), .Y(n7325) );
  MUX2X1 U10614 ( .B(n7324), .A(n7309), .S(N17), .Y(n8318) );
  MUX2X1 U10615 ( .B(\RF[30][32] ), .A(\RF[31][32] ), .S(n8414), .Y(n7329) );
  MUX2X1 U10616 ( .B(\RF[28][32] ), .A(\RF[29][32] ), .S(n8414), .Y(n7328) );
  MUX2X1 U10617 ( .B(\RF[26][32] ), .A(\RF[27][32] ), .S(n8414), .Y(n7332) );
  MUX2X1 U10618 ( .B(\RF[24][32] ), .A(\RF[25][32] ), .S(n8414), .Y(n7331) );
  MUX2X1 U10619 ( .B(n7330), .A(n7327), .S(n8526), .Y(n7341) );
  MUX2X1 U10620 ( .B(\RF[22][32] ), .A(\RF[23][32] ), .S(n8414), .Y(n7335) );
  MUX2X1 U10621 ( .B(\RF[20][32] ), .A(\RF[21][32] ), .S(n8414), .Y(n7334) );
  MUX2X1 U10622 ( .B(\RF[18][32] ), .A(\RF[19][32] ), .S(n8414), .Y(n7338) );
  MUX2X1 U10623 ( .B(\RF[16][32] ), .A(\RF[17][32] ), .S(n8414), .Y(n7337) );
  MUX2X1 U10624 ( .B(n7336), .A(n7333), .S(n8526), .Y(n7340) );
  MUX2X1 U10625 ( .B(\RF[14][32] ), .A(\RF[15][32] ), .S(n8415), .Y(n7344) );
  MUX2X1 U10626 ( .B(\RF[12][32] ), .A(\RF[13][32] ), .S(n8415), .Y(n7343) );
  MUX2X1 U10627 ( .B(\RF[10][32] ), .A(\RF[11][32] ), .S(n8415), .Y(n7347) );
  MUX2X1 U10628 ( .B(\RF[8][32] ), .A(\RF[9][32] ), .S(n8415), .Y(n7346) );
  MUX2X1 U10629 ( .B(n7345), .A(n7342), .S(n8526), .Y(n7356) );
  MUX2X1 U10630 ( .B(\RF[6][32] ), .A(\RF[7][32] ), .S(n8415), .Y(n7350) );
  MUX2X1 U10631 ( .B(\RF[4][32] ), .A(\RF[5][32] ), .S(n8415), .Y(n7349) );
  MUX2X1 U10632 ( .B(\RF[2][32] ), .A(\RF[3][32] ), .S(n8415), .Y(n7353) );
  MUX2X1 U10633 ( .B(\RF[0][32] ), .A(\RF[1][32] ), .S(n8415), .Y(n7352) );
  MUX2X1 U10634 ( .B(n7351), .A(n7348), .S(n8526), .Y(n7355) );
  MUX2X1 U10635 ( .B(n7354), .A(n7339), .S(N17), .Y(n8319) );
  MUX2X1 U10636 ( .B(\RF[30][33] ), .A(\RF[31][33] ), .S(n8415), .Y(n7359) );
  MUX2X1 U10637 ( .B(\RF[28][33] ), .A(\RF[29][33] ), .S(n8415), .Y(n7358) );
  MUX2X1 U10638 ( .B(\RF[26][33] ), .A(\RF[27][33] ), .S(n8415), .Y(n7362) );
  MUX2X1 U10639 ( .B(\RF[24][33] ), .A(\RF[25][33] ), .S(n8415), .Y(n7361) );
  MUX2X1 U10640 ( .B(n7360), .A(n7357), .S(n8526), .Y(n7371) );
  MUX2X1 U10641 ( .B(\RF[22][33] ), .A(\RF[23][33] ), .S(n8416), .Y(n7365) );
  MUX2X1 U10642 ( .B(\RF[20][33] ), .A(\RF[21][33] ), .S(n8416), .Y(n7364) );
  MUX2X1 U10643 ( .B(\RF[18][33] ), .A(\RF[19][33] ), .S(n8416), .Y(n7368) );
  MUX2X1 U10644 ( .B(\RF[16][33] ), .A(\RF[17][33] ), .S(n8416), .Y(n7367) );
  MUX2X1 U10645 ( .B(n7366), .A(n7363), .S(n8526), .Y(n7370) );
  MUX2X1 U10646 ( .B(\RF[14][33] ), .A(\RF[15][33] ), .S(n8416), .Y(n7374) );
  MUX2X1 U10647 ( .B(\RF[12][33] ), .A(\RF[13][33] ), .S(n8416), .Y(n7373) );
  MUX2X1 U10648 ( .B(\RF[10][33] ), .A(\RF[11][33] ), .S(n8416), .Y(n7377) );
  MUX2X1 U10649 ( .B(\RF[8][33] ), .A(\RF[9][33] ), .S(n8416), .Y(n7376) );
  MUX2X1 U10650 ( .B(n7375), .A(n7372), .S(n8526), .Y(n7386) );
  MUX2X1 U10651 ( .B(\RF[6][33] ), .A(\RF[7][33] ), .S(n8416), .Y(n7380) );
  MUX2X1 U10652 ( .B(\RF[4][33] ), .A(\RF[5][33] ), .S(n8416), .Y(n7379) );
  MUX2X1 U10653 ( .B(\RF[2][33] ), .A(\RF[3][33] ), .S(n8416), .Y(n7383) );
  MUX2X1 U10654 ( .B(\RF[0][33] ), .A(\RF[1][33] ), .S(n8416), .Y(n7382) );
  MUX2X1 U10655 ( .B(n7381), .A(n7378), .S(n8526), .Y(n7385) );
  MUX2X1 U10656 ( .B(n7384), .A(n7369), .S(N17), .Y(n8320) );
  MUX2X1 U10657 ( .B(\RF[30][34] ), .A(\RF[31][34] ), .S(n8417), .Y(n7389) );
  MUX2X1 U10658 ( .B(\RF[28][34] ), .A(\RF[29][34] ), .S(n8417), .Y(n7388) );
  MUX2X1 U10659 ( .B(\RF[26][34] ), .A(\RF[27][34] ), .S(n8417), .Y(n7392) );
  MUX2X1 U10660 ( .B(\RF[24][34] ), .A(\RF[25][34] ), .S(n8417), .Y(n7391) );
  MUX2X1 U10661 ( .B(n7390), .A(n7387), .S(n8527), .Y(n7401) );
  MUX2X1 U10662 ( .B(\RF[22][34] ), .A(\RF[23][34] ), .S(n8417), .Y(n7395) );
  MUX2X1 U10663 ( .B(\RF[20][34] ), .A(\RF[21][34] ), .S(n8417), .Y(n7394) );
  MUX2X1 U10664 ( .B(\RF[18][34] ), .A(\RF[19][34] ), .S(n8417), .Y(n7398) );
  MUX2X1 U10665 ( .B(\RF[16][34] ), .A(\RF[17][34] ), .S(n8417), .Y(n7397) );
  MUX2X1 U10666 ( .B(n7396), .A(n7393), .S(n8527), .Y(n7400) );
  MUX2X1 U10667 ( .B(\RF[14][34] ), .A(\RF[15][34] ), .S(n8417), .Y(n7404) );
  MUX2X1 U10668 ( .B(\RF[12][34] ), .A(\RF[13][34] ), .S(n8417), .Y(n7403) );
  MUX2X1 U10669 ( .B(\RF[10][34] ), .A(\RF[11][34] ), .S(n8417), .Y(n7407) );
  MUX2X1 U10670 ( .B(\RF[8][34] ), .A(\RF[9][34] ), .S(n8417), .Y(n7406) );
  MUX2X1 U10671 ( .B(n7405), .A(n7402), .S(n8527), .Y(n7416) );
  MUX2X1 U10672 ( .B(\RF[6][34] ), .A(\RF[7][34] ), .S(n8418), .Y(n7410) );
  MUX2X1 U10673 ( .B(\RF[4][34] ), .A(\RF[5][34] ), .S(n8418), .Y(n7409) );
  MUX2X1 U10674 ( .B(\RF[2][34] ), .A(\RF[3][34] ), .S(n8418), .Y(n7413) );
  MUX2X1 U10675 ( .B(\RF[0][34] ), .A(\RF[1][34] ), .S(n8418), .Y(n7412) );
  MUX2X1 U10676 ( .B(n7411), .A(n7408), .S(n8527), .Y(n7415) );
  MUX2X1 U10677 ( .B(n7414), .A(n7399), .S(N17), .Y(n8321) );
  MUX2X1 U10678 ( .B(\RF[30][35] ), .A(\RF[31][35] ), .S(n8418), .Y(n7419) );
  MUX2X1 U10679 ( .B(\RF[28][35] ), .A(\RF[29][35] ), .S(n8418), .Y(n7418) );
  MUX2X1 U10680 ( .B(\RF[26][35] ), .A(\RF[27][35] ), .S(n8418), .Y(n7422) );
  MUX2X1 U10681 ( .B(\RF[24][35] ), .A(\RF[25][35] ), .S(n8418), .Y(n7421) );
  MUX2X1 U10682 ( .B(n7420), .A(n7417), .S(n8527), .Y(n7431) );
  MUX2X1 U10683 ( .B(\RF[22][35] ), .A(\RF[23][35] ), .S(n8418), .Y(n7425) );
  MUX2X1 U10684 ( .B(\RF[20][35] ), .A(\RF[21][35] ), .S(n8418), .Y(n7424) );
  MUX2X1 U10685 ( .B(\RF[18][35] ), .A(\RF[19][35] ), .S(n8418), .Y(n7428) );
  MUX2X1 U10686 ( .B(\RF[16][35] ), .A(\RF[17][35] ), .S(n8418), .Y(n7427) );
  MUX2X1 U10687 ( .B(n7426), .A(n7423), .S(n8527), .Y(n7430) );
  MUX2X1 U10688 ( .B(\RF[14][35] ), .A(\RF[15][35] ), .S(n8419), .Y(n7434) );
  MUX2X1 U10689 ( .B(\RF[12][35] ), .A(\RF[13][35] ), .S(n8419), .Y(n7433) );
  MUX2X1 U10690 ( .B(\RF[10][35] ), .A(\RF[11][35] ), .S(n8419), .Y(n7437) );
  MUX2X1 U10691 ( .B(\RF[8][35] ), .A(\RF[9][35] ), .S(n8419), .Y(n7436) );
  MUX2X1 U10692 ( .B(n7435), .A(n7432), .S(n8527), .Y(n7446) );
  MUX2X1 U10693 ( .B(\RF[6][35] ), .A(\RF[7][35] ), .S(n8419), .Y(n7440) );
  MUX2X1 U10694 ( .B(\RF[4][35] ), .A(\RF[5][35] ), .S(n8419), .Y(n7439) );
  MUX2X1 U10695 ( .B(\RF[2][35] ), .A(\RF[3][35] ), .S(n8419), .Y(n7443) );
  MUX2X1 U10696 ( .B(\RF[0][35] ), .A(\RF[1][35] ), .S(n8419), .Y(n7442) );
  MUX2X1 U10697 ( .B(n7441), .A(n7438), .S(n8527), .Y(n7445) );
  MUX2X1 U10698 ( .B(n7444), .A(n7429), .S(N17), .Y(n8322) );
  MUX2X1 U10699 ( .B(\RF[30][36] ), .A(\RF[31][36] ), .S(n8419), .Y(n7449) );
  MUX2X1 U10700 ( .B(\RF[28][36] ), .A(\RF[29][36] ), .S(n8419), .Y(n7448) );
  MUX2X1 U10701 ( .B(\RF[26][36] ), .A(\RF[27][36] ), .S(n8419), .Y(n7452) );
  MUX2X1 U10702 ( .B(\RF[24][36] ), .A(\RF[25][36] ), .S(n8419), .Y(n7451) );
  MUX2X1 U10703 ( .B(n7450), .A(n7447), .S(n8527), .Y(n7461) );
  MUX2X1 U10704 ( .B(\RF[22][36] ), .A(\RF[23][36] ), .S(n8420), .Y(n7455) );
  MUX2X1 U10705 ( .B(\RF[20][36] ), .A(\RF[21][36] ), .S(n8420), .Y(n7454) );
  MUX2X1 U10706 ( .B(\RF[18][36] ), .A(\RF[19][36] ), .S(n8420), .Y(n7458) );
  MUX2X1 U10707 ( .B(\RF[16][36] ), .A(\RF[17][36] ), .S(n8420), .Y(n7457) );
  MUX2X1 U10708 ( .B(n7456), .A(n7453), .S(n8527), .Y(n7460) );
  MUX2X1 U10709 ( .B(\RF[14][36] ), .A(\RF[15][36] ), .S(n8420), .Y(n7464) );
  MUX2X1 U10710 ( .B(\RF[12][36] ), .A(\RF[13][36] ), .S(n8420), .Y(n7463) );
  MUX2X1 U10711 ( .B(\RF[10][36] ), .A(\RF[11][36] ), .S(n8420), .Y(n7467) );
  MUX2X1 U10712 ( .B(\RF[8][36] ), .A(\RF[9][36] ), .S(n8420), .Y(n7466) );
  MUX2X1 U10713 ( .B(n7465), .A(n7462), .S(n8527), .Y(n7476) );
  MUX2X1 U10714 ( .B(\RF[6][36] ), .A(\RF[7][36] ), .S(n8420), .Y(n7470) );
  MUX2X1 U10715 ( .B(\RF[4][36] ), .A(\RF[5][36] ), .S(n8420), .Y(n7469) );
  MUX2X1 U10716 ( .B(\RF[2][36] ), .A(\RF[3][36] ), .S(n8420), .Y(n7473) );
  MUX2X1 U10717 ( .B(\RF[0][36] ), .A(\RF[1][36] ), .S(n8420), .Y(n7472) );
  MUX2X1 U10718 ( .B(n7471), .A(n7468), .S(n8527), .Y(n7475) );
  MUX2X1 U10719 ( .B(n7474), .A(n7459), .S(N17), .Y(n8323) );
  MUX2X1 U10720 ( .B(\RF[30][37] ), .A(\RF[31][37] ), .S(n8421), .Y(n7479) );
  MUX2X1 U10721 ( .B(\RF[28][37] ), .A(\RF[29][37] ), .S(n8421), .Y(n7478) );
  MUX2X1 U10722 ( .B(\RF[26][37] ), .A(\RF[27][37] ), .S(n8421), .Y(n7482) );
  MUX2X1 U10723 ( .B(\RF[24][37] ), .A(\RF[25][37] ), .S(n8421), .Y(n7481) );
  MUX2X1 U10724 ( .B(n7480), .A(n7477), .S(n8528), .Y(n7491) );
  MUX2X1 U10725 ( .B(\RF[22][37] ), .A(\RF[23][37] ), .S(n8421), .Y(n7485) );
  MUX2X1 U10726 ( .B(\RF[20][37] ), .A(\RF[21][37] ), .S(n8421), .Y(n7484) );
  MUX2X1 U10727 ( .B(\RF[18][37] ), .A(\RF[19][37] ), .S(n8421), .Y(n7488) );
  MUX2X1 U10728 ( .B(\RF[16][37] ), .A(\RF[17][37] ), .S(n8421), .Y(n7487) );
  MUX2X1 U10729 ( .B(n7486), .A(n7483), .S(n8528), .Y(n7490) );
  MUX2X1 U10730 ( .B(\RF[14][37] ), .A(\RF[15][37] ), .S(n8421), .Y(n7494) );
  MUX2X1 U10731 ( .B(\RF[12][37] ), .A(\RF[13][37] ), .S(n8421), .Y(n7493) );
  MUX2X1 U10732 ( .B(\RF[10][37] ), .A(\RF[11][37] ), .S(n8421), .Y(n7497) );
  MUX2X1 U10733 ( .B(\RF[8][37] ), .A(\RF[9][37] ), .S(n8421), .Y(n7496) );
  MUX2X1 U10734 ( .B(n7495), .A(n7492), .S(n8528), .Y(n7506) );
  MUX2X1 U10735 ( .B(\RF[6][37] ), .A(\RF[7][37] ), .S(n8422), .Y(n7500) );
  MUX2X1 U10736 ( .B(\RF[4][37] ), .A(\RF[5][37] ), .S(n8422), .Y(n7499) );
  MUX2X1 U10737 ( .B(\RF[2][37] ), .A(\RF[3][37] ), .S(n8422), .Y(n7503) );
  MUX2X1 U10738 ( .B(\RF[0][37] ), .A(\RF[1][37] ), .S(n8422), .Y(n7502) );
  MUX2X1 U10739 ( .B(n7501), .A(n7498), .S(n8528), .Y(n7505) );
  MUX2X1 U10740 ( .B(n7504), .A(n7489), .S(N17), .Y(n8324) );
  MUX2X1 U10741 ( .B(\RF[30][38] ), .A(\RF[31][38] ), .S(n8422), .Y(n7509) );
  MUX2X1 U10742 ( .B(\RF[28][38] ), .A(\RF[29][38] ), .S(n8422), .Y(n7508) );
  MUX2X1 U10743 ( .B(\RF[26][38] ), .A(\RF[27][38] ), .S(n8422), .Y(n7512) );
  MUX2X1 U10744 ( .B(\RF[24][38] ), .A(\RF[25][38] ), .S(n8422), .Y(n7511) );
  MUX2X1 U10745 ( .B(n7510), .A(n7507), .S(n8528), .Y(n7521) );
  MUX2X1 U10746 ( .B(\RF[22][38] ), .A(\RF[23][38] ), .S(n8422), .Y(n7515) );
  MUX2X1 U10747 ( .B(\RF[20][38] ), .A(\RF[21][38] ), .S(n8422), .Y(n7514) );
  MUX2X1 U10748 ( .B(\RF[18][38] ), .A(\RF[19][38] ), .S(n8422), .Y(n7518) );
  MUX2X1 U10749 ( .B(\RF[16][38] ), .A(\RF[17][38] ), .S(n8422), .Y(n7517) );
  MUX2X1 U10750 ( .B(n7516), .A(n7513), .S(n8528), .Y(n7520) );
  MUX2X1 U10751 ( .B(\RF[14][38] ), .A(\RF[15][38] ), .S(n8423), .Y(n7524) );
  MUX2X1 U10752 ( .B(\RF[12][38] ), .A(\RF[13][38] ), .S(n8423), .Y(n7523) );
  MUX2X1 U10753 ( .B(\RF[10][38] ), .A(\RF[11][38] ), .S(n8423), .Y(n7527) );
  MUX2X1 U10754 ( .B(\RF[8][38] ), .A(\RF[9][38] ), .S(n8423), .Y(n7526) );
  MUX2X1 U10755 ( .B(n7525), .A(n7522), .S(n8528), .Y(n7536) );
  MUX2X1 U10756 ( .B(\RF[6][38] ), .A(\RF[7][38] ), .S(n8423), .Y(n7530) );
  MUX2X1 U10757 ( .B(\RF[4][38] ), .A(\RF[5][38] ), .S(n8423), .Y(n7529) );
  MUX2X1 U10758 ( .B(\RF[2][38] ), .A(\RF[3][38] ), .S(n8423), .Y(n7533) );
  MUX2X1 U10759 ( .B(\RF[0][38] ), .A(\RF[1][38] ), .S(n8423), .Y(n7532) );
  MUX2X1 U10760 ( .B(n7531), .A(n7528), .S(n8528), .Y(n7535) );
  MUX2X1 U10761 ( .B(n7534), .A(n7519), .S(N17), .Y(n8325) );
  MUX2X1 U10762 ( .B(\RF[30][39] ), .A(\RF[31][39] ), .S(n8423), .Y(n7539) );
  MUX2X1 U10763 ( .B(\RF[28][39] ), .A(\RF[29][39] ), .S(n8423), .Y(n7538) );
  MUX2X1 U10764 ( .B(\RF[26][39] ), .A(\RF[27][39] ), .S(n8423), .Y(n7542) );
  MUX2X1 U10765 ( .B(\RF[24][39] ), .A(\RF[25][39] ), .S(n8423), .Y(n7541) );
  MUX2X1 U10766 ( .B(n7540), .A(n7537), .S(n8528), .Y(n7551) );
  MUX2X1 U10767 ( .B(\RF[22][39] ), .A(\RF[23][39] ), .S(n8424), .Y(n7545) );
  MUX2X1 U10768 ( .B(\RF[20][39] ), .A(\RF[21][39] ), .S(n8424), .Y(n7544) );
  MUX2X1 U10769 ( .B(\RF[18][39] ), .A(\RF[19][39] ), .S(n8424), .Y(n7548) );
  MUX2X1 U10770 ( .B(\RF[16][39] ), .A(\RF[17][39] ), .S(n8424), .Y(n7547) );
  MUX2X1 U10771 ( .B(n7546), .A(n7543), .S(n8528), .Y(n7550) );
  MUX2X1 U10772 ( .B(\RF[14][39] ), .A(\RF[15][39] ), .S(n8424), .Y(n7554) );
  MUX2X1 U10773 ( .B(\RF[12][39] ), .A(\RF[13][39] ), .S(n8424), .Y(n7553) );
  MUX2X1 U10774 ( .B(\RF[10][39] ), .A(\RF[11][39] ), .S(n8424), .Y(n7557) );
  MUX2X1 U10775 ( .B(\RF[8][39] ), .A(\RF[9][39] ), .S(n8424), .Y(n7556) );
  MUX2X1 U10776 ( .B(n7555), .A(n7552), .S(n8528), .Y(n7566) );
  MUX2X1 U10777 ( .B(\RF[6][39] ), .A(\RF[7][39] ), .S(n8424), .Y(n7560) );
  MUX2X1 U10778 ( .B(\RF[4][39] ), .A(\RF[5][39] ), .S(n8424), .Y(n7559) );
  MUX2X1 U10779 ( .B(\RF[2][39] ), .A(\RF[3][39] ), .S(n8424), .Y(n7563) );
  MUX2X1 U10780 ( .B(\RF[0][39] ), .A(\RF[1][39] ), .S(n8424), .Y(n7562) );
  MUX2X1 U10781 ( .B(n7561), .A(n7558), .S(n8528), .Y(n7565) );
  MUX2X1 U10782 ( .B(n7564), .A(n7549), .S(N17), .Y(n8326) );
  MUX2X1 U10783 ( .B(\RF[30][40] ), .A(\RF[31][40] ), .S(n8425), .Y(n7569) );
  MUX2X1 U10784 ( .B(\RF[28][40] ), .A(\RF[29][40] ), .S(n8425), .Y(n7568) );
  MUX2X1 U10785 ( .B(\RF[26][40] ), .A(\RF[27][40] ), .S(n8425), .Y(n7572) );
  MUX2X1 U10786 ( .B(\RF[24][40] ), .A(\RF[25][40] ), .S(n8425), .Y(n7571) );
  MUX2X1 U10787 ( .B(n7570), .A(n7567), .S(n8529), .Y(n7581) );
  MUX2X1 U10788 ( .B(\RF[22][40] ), .A(\RF[23][40] ), .S(n8425), .Y(n7575) );
  MUX2X1 U10789 ( .B(\RF[20][40] ), .A(\RF[21][40] ), .S(n8425), .Y(n7574) );
  MUX2X1 U10790 ( .B(\RF[18][40] ), .A(\RF[19][40] ), .S(n8425), .Y(n7578) );
  MUX2X1 U10791 ( .B(\RF[16][40] ), .A(\RF[17][40] ), .S(n8425), .Y(n7577) );
  MUX2X1 U10792 ( .B(n7576), .A(n7573), .S(n8529), .Y(n7580) );
  MUX2X1 U10793 ( .B(\RF[14][40] ), .A(\RF[15][40] ), .S(n8425), .Y(n7584) );
  MUX2X1 U10794 ( .B(\RF[12][40] ), .A(\RF[13][40] ), .S(n8425), .Y(n7583) );
  MUX2X1 U10795 ( .B(\RF[10][40] ), .A(\RF[11][40] ), .S(n8425), .Y(n7587) );
  MUX2X1 U10796 ( .B(\RF[8][40] ), .A(\RF[9][40] ), .S(n8425), .Y(n7586) );
  MUX2X1 U10797 ( .B(n7585), .A(n7582), .S(n8529), .Y(n7596) );
  MUX2X1 U10798 ( .B(\RF[6][40] ), .A(\RF[7][40] ), .S(n8426), .Y(n7590) );
  MUX2X1 U10799 ( .B(\RF[4][40] ), .A(\RF[5][40] ), .S(n8426), .Y(n7589) );
  MUX2X1 U10800 ( .B(\RF[2][40] ), .A(\RF[3][40] ), .S(n8426), .Y(n7593) );
  MUX2X1 U10801 ( .B(\RF[0][40] ), .A(\RF[1][40] ), .S(n8426), .Y(n7592) );
  MUX2X1 U10802 ( .B(n7591), .A(n7588), .S(n8529), .Y(n7595) );
  MUX2X1 U10803 ( .B(n7594), .A(n7579), .S(N17), .Y(n8327) );
  MUX2X1 U10804 ( .B(\RF[30][41] ), .A(\RF[31][41] ), .S(n8426), .Y(n7599) );
  MUX2X1 U10805 ( .B(\RF[28][41] ), .A(\RF[29][41] ), .S(n8426), .Y(n7598) );
  MUX2X1 U10806 ( .B(\RF[26][41] ), .A(\RF[27][41] ), .S(n8426), .Y(n7602) );
  MUX2X1 U10807 ( .B(\RF[24][41] ), .A(\RF[25][41] ), .S(n8426), .Y(n7601) );
  MUX2X1 U10808 ( .B(n7600), .A(n7597), .S(n8529), .Y(n7611) );
  MUX2X1 U10809 ( .B(\RF[22][41] ), .A(\RF[23][41] ), .S(n8426), .Y(n7605) );
  MUX2X1 U10810 ( .B(\RF[20][41] ), .A(\RF[21][41] ), .S(n8426), .Y(n7604) );
  MUX2X1 U10811 ( .B(\RF[18][41] ), .A(\RF[19][41] ), .S(n8426), .Y(n7608) );
  MUX2X1 U10812 ( .B(\RF[16][41] ), .A(\RF[17][41] ), .S(n8426), .Y(n7607) );
  MUX2X1 U10813 ( .B(n7606), .A(n7603), .S(n8529), .Y(n7610) );
  MUX2X1 U10814 ( .B(\RF[14][41] ), .A(\RF[15][41] ), .S(n8427), .Y(n7614) );
  MUX2X1 U10815 ( .B(\RF[12][41] ), .A(\RF[13][41] ), .S(n8427), .Y(n7613) );
  MUX2X1 U10816 ( .B(\RF[10][41] ), .A(\RF[11][41] ), .S(n8427), .Y(n7617) );
  MUX2X1 U10817 ( .B(\RF[8][41] ), .A(\RF[9][41] ), .S(n8427), .Y(n7616) );
  MUX2X1 U10818 ( .B(n7615), .A(n7612), .S(n8529), .Y(n7626) );
  MUX2X1 U10819 ( .B(\RF[6][41] ), .A(\RF[7][41] ), .S(n8427), .Y(n7620) );
  MUX2X1 U10820 ( .B(\RF[4][41] ), .A(\RF[5][41] ), .S(n8427), .Y(n7619) );
  MUX2X1 U10821 ( .B(\RF[2][41] ), .A(\RF[3][41] ), .S(n8427), .Y(n7623) );
  MUX2X1 U10822 ( .B(\RF[0][41] ), .A(\RF[1][41] ), .S(n8427), .Y(n7622) );
  MUX2X1 U10823 ( .B(n7621), .A(n7618), .S(n8529), .Y(n7625) );
  MUX2X1 U10824 ( .B(n7624), .A(n7609), .S(N17), .Y(n8328) );
  MUX2X1 U10825 ( .B(\RF[30][42] ), .A(\RF[31][42] ), .S(n8427), .Y(n7629) );
  MUX2X1 U10826 ( .B(\RF[28][42] ), .A(\RF[29][42] ), .S(n8427), .Y(n7628) );
  MUX2X1 U10827 ( .B(\RF[26][42] ), .A(\RF[27][42] ), .S(n8427), .Y(n7632) );
  MUX2X1 U10828 ( .B(\RF[24][42] ), .A(\RF[25][42] ), .S(n8427), .Y(n7631) );
  MUX2X1 U10829 ( .B(n7630), .A(n7627), .S(n8529), .Y(n7641) );
  MUX2X1 U10830 ( .B(\RF[22][42] ), .A(\RF[23][42] ), .S(n8428), .Y(n7635) );
  MUX2X1 U10831 ( .B(\RF[20][42] ), .A(\RF[21][42] ), .S(n8428), .Y(n7634) );
  MUX2X1 U10832 ( .B(\RF[18][42] ), .A(\RF[19][42] ), .S(n8428), .Y(n7638) );
  MUX2X1 U10833 ( .B(\RF[16][42] ), .A(\RF[17][42] ), .S(n8428), .Y(n7637) );
  MUX2X1 U10834 ( .B(n7636), .A(n7633), .S(n8529), .Y(n7640) );
  MUX2X1 U10835 ( .B(\RF[14][42] ), .A(\RF[15][42] ), .S(n8428), .Y(n7644) );
  MUX2X1 U10836 ( .B(\RF[12][42] ), .A(\RF[13][42] ), .S(n8428), .Y(n7643) );
  MUX2X1 U10837 ( .B(\RF[10][42] ), .A(\RF[11][42] ), .S(n8428), .Y(n7647) );
  MUX2X1 U10838 ( .B(\RF[8][42] ), .A(\RF[9][42] ), .S(n8428), .Y(n7646) );
  MUX2X1 U10839 ( .B(n7645), .A(n7642), .S(n8529), .Y(n7656) );
  MUX2X1 U10840 ( .B(\RF[6][42] ), .A(\RF[7][42] ), .S(n8428), .Y(n7650) );
  MUX2X1 U10841 ( .B(\RF[4][42] ), .A(\RF[5][42] ), .S(n8428), .Y(n7649) );
  MUX2X1 U10842 ( .B(\RF[2][42] ), .A(\RF[3][42] ), .S(n8428), .Y(n7653) );
  MUX2X1 U10843 ( .B(\RF[0][42] ), .A(\RF[1][42] ), .S(n8428), .Y(n7652) );
  MUX2X1 U10844 ( .B(n7651), .A(n7648), .S(n8529), .Y(n7655) );
  MUX2X1 U10845 ( .B(n7654), .A(n7639), .S(N17), .Y(n8329) );
  MUX2X1 U10846 ( .B(\RF[30][43] ), .A(\RF[31][43] ), .S(n8429), .Y(n7659) );
  MUX2X1 U10847 ( .B(\RF[28][43] ), .A(\RF[29][43] ), .S(n8429), .Y(n7658) );
  MUX2X1 U10848 ( .B(\RF[26][43] ), .A(\RF[27][43] ), .S(n8429), .Y(n7662) );
  MUX2X1 U10849 ( .B(\RF[24][43] ), .A(\RF[25][43] ), .S(n8429), .Y(n7661) );
  MUX2X1 U10850 ( .B(n7660), .A(n7657), .S(n8530), .Y(n7671) );
  MUX2X1 U10851 ( .B(\RF[22][43] ), .A(\RF[23][43] ), .S(n8429), .Y(n7665) );
  MUX2X1 U10852 ( .B(\RF[20][43] ), .A(\RF[21][43] ), .S(n8429), .Y(n7664) );
  MUX2X1 U10853 ( .B(\RF[18][43] ), .A(\RF[19][43] ), .S(n8429), .Y(n7668) );
  MUX2X1 U10854 ( .B(\RF[16][43] ), .A(\RF[17][43] ), .S(n8429), .Y(n7667) );
  MUX2X1 U10855 ( .B(n7666), .A(n7663), .S(n8530), .Y(n7670) );
  MUX2X1 U10856 ( .B(\RF[14][43] ), .A(\RF[15][43] ), .S(n8429), .Y(n7674) );
  MUX2X1 U10857 ( .B(\RF[12][43] ), .A(\RF[13][43] ), .S(n8429), .Y(n7673) );
  MUX2X1 U10858 ( .B(\RF[10][43] ), .A(\RF[11][43] ), .S(n8429), .Y(n7677) );
  MUX2X1 U10859 ( .B(\RF[8][43] ), .A(\RF[9][43] ), .S(n8429), .Y(n7676) );
  MUX2X1 U10860 ( .B(n7675), .A(n7672), .S(n8530), .Y(n7686) );
  MUX2X1 U10861 ( .B(\RF[6][43] ), .A(\RF[7][43] ), .S(n8430), .Y(n7680) );
  MUX2X1 U10862 ( .B(\RF[4][43] ), .A(\RF[5][43] ), .S(n8430), .Y(n7679) );
  MUX2X1 U10863 ( .B(\RF[2][43] ), .A(\RF[3][43] ), .S(n8430), .Y(n7683) );
  MUX2X1 U10864 ( .B(\RF[0][43] ), .A(\RF[1][43] ), .S(n8430), .Y(n7682) );
  MUX2X1 U10865 ( .B(n7681), .A(n7678), .S(n8530), .Y(n7685) );
  MUX2X1 U10866 ( .B(n7684), .A(n7669), .S(N17), .Y(n8330) );
  MUX2X1 U10867 ( .B(\RF[30][44] ), .A(\RF[31][44] ), .S(n8430), .Y(n7689) );
  MUX2X1 U10868 ( .B(\RF[28][44] ), .A(\RF[29][44] ), .S(n8430), .Y(n7688) );
  MUX2X1 U10869 ( .B(\RF[26][44] ), .A(\RF[27][44] ), .S(n8430), .Y(n7692) );
  MUX2X1 U10870 ( .B(\RF[24][44] ), .A(\RF[25][44] ), .S(n8430), .Y(n7691) );
  MUX2X1 U10871 ( .B(n7690), .A(n7687), .S(n8530), .Y(n7701) );
  MUX2X1 U10872 ( .B(\RF[22][44] ), .A(\RF[23][44] ), .S(n8430), .Y(n7695) );
  MUX2X1 U10873 ( .B(\RF[20][44] ), .A(\RF[21][44] ), .S(n8430), .Y(n7694) );
  MUX2X1 U10874 ( .B(\RF[18][44] ), .A(\RF[19][44] ), .S(n8430), .Y(n7698) );
  MUX2X1 U10875 ( .B(\RF[16][44] ), .A(\RF[17][44] ), .S(n8430), .Y(n7697) );
  MUX2X1 U10876 ( .B(n7696), .A(n7693), .S(n8530), .Y(n7700) );
  MUX2X1 U10877 ( .B(\RF[14][44] ), .A(\RF[15][44] ), .S(n8431), .Y(n7704) );
  MUX2X1 U10878 ( .B(\RF[12][44] ), .A(\RF[13][44] ), .S(n8431), .Y(n7703) );
  MUX2X1 U10879 ( .B(\RF[10][44] ), .A(\RF[11][44] ), .S(n8431), .Y(n7707) );
  MUX2X1 U10880 ( .B(\RF[8][44] ), .A(\RF[9][44] ), .S(n8431), .Y(n7706) );
  MUX2X1 U10881 ( .B(n7705), .A(n7702), .S(n8530), .Y(n7716) );
  MUX2X1 U10882 ( .B(\RF[6][44] ), .A(\RF[7][44] ), .S(n8431), .Y(n7710) );
  MUX2X1 U10883 ( .B(\RF[4][44] ), .A(\RF[5][44] ), .S(n8431), .Y(n7709) );
  MUX2X1 U10884 ( .B(\RF[2][44] ), .A(\RF[3][44] ), .S(n8431), .Y(n7713) );
  MUX2X1 U10885 ( .B(\RF[0][44] ), .A(\RF[1][44] ), .S(n8431), .Y(n7712) );
  MUX2X1 U10886 ( .B(n7711), .A(n7708), .S(n8530), .Y(n7715) );
  MUX2X1 U10887 ( .B(n7714), .A(n7699), .S(N17), .Y(n8331) );
  MUX2X1 U10888 ( .B(\RF[30][45] ), .A(\RF[31][45] ), .S(n8431), .Y(n7719) );
  MUX2X1 U10889 ( .B(\RF[28][45] ), .A(\RF[29][45] ), .S(n8431), .Y(n7718) );
  MUX2X1 U10890 ( .B(\RF[26][45] ), .A(\RF[27][45] ), .S(n8431), .Y(n7722) );
  MUX2X1 U10891 ( .B(\RF[24][45] ), .A(\RF[25][45] ), .S(n8431), .Y(n7721) );
  MUX2X1 U10892 ( .B(n7720), .A(n7717), .S(n8530), .Y(n7731) );
  MUX2X1 U10893 ( .B(\RF[22][45] ), .A(\RF[23][45] ), .S(n8432), .Y(n7725) );
  MUX2X1 U10894 ( .B(\RF[20][45] ), .A(\RF[21][45] ), .S(n8432), .Y(n7724) );
  MUX2X1 U10895 ( .B(\RF[18][45] ), .A(\RF[19][45] ), .S(n8432), .Y(n7728) );
  MUX2X1 U10896 ( .B(\RF[16][45] ), .A(\RF[17][45] ), .S(n8432), .Y(n7727) );
  MUX2X1 U10897 ( .B(n7726), .A(n7723), .S(n8530), .Y(n7730) );
  MUX2X1 U10898 ( .B(\RF[14][45] ), .A(\RF[15][45] ), .S(n8432), .Y(n7734) );
  MUX2X1 U10899 ( .B(\RF[12][45] ), .A(\RF[13][45] ), .S(n8432), .Y(n7733) );
  MUX2X1 U10900 ( .B(\RF[10][45] ), .A(\RF[11][45] ), .S(n8432), .Y(n7737) );
  MUX2X1 U10901 ( .B(\RF[8][45] ), .A(\RF[9][45] ), .S(n8432), .Y(n7736) );
  MUX2X1 U10902 ( .B(n7735), .A(n7732), .S(n8530), .Y(n7746) );
  MUX2X1 U10903 ( .B(\RF[6][45] ), .A(\RF[7][45] ), .S(n8432), .Y(n7740) );
  MUX2X1 U10904 ( .B(\RF[4][45] ), .A(\RF[5][45] ), .S(n8432), .Y(n7739) );
  MUX2X1 U10905 ( .B(\RF[2][45] ), .A(\RF[3][45] ), .S(n8432), .Y(n7743) );
  MUX2X1 U10906 ( .B(\RF[0][45] ), .A(\RF[1][45] ), .S(n8432), .Y(n7742) );
  MUX2X1 U10907 ( .B(n7741), .A(n7738), .S(n8530), .Y(n7745) );
  MUX2X1 U10908 ( .B(n7744), .A(n7729), .S(N17), .Y(n8332) );
  MUX2X1 U10909 ( .B(\RF[30][46] ), .A(\RF[31][46] ), .S(n8433), .Y(n7749) );
  MUX2X1 U10910 ( .B(\RF[28][46] ), .A(\RF[29][46] ), .S(n8433), .Y(n7748) );
  MUX2X1 U10911 ( .B(\RF[26][46] ), .A(\RF[27][46] ), .S(n8433), .Y(n7752) );
  MUX2X1 U10912 ( .B(\RF[24][46] ), .A(\RF[25][46] ), .S(n8433), .Y(n7751) );
  MUX2X1 U10913 ( .B(n7750), .A(n7747), .S(n8531), .Y(n7761) );
  MUX2X1 U10914 ( .B(\RF[22][46] ), .A(\RF[23][46] ), .S(n8433), .Y(n7755) );
  MUX2X1 U10915 ( .B(\RF[20][46] ), .A(\RF[21][46] ), .S(n8433), .Y(n7754) );
  MUX2X1 U10916 ( .B(\RF[18][46] ), .A(\RF[19][46] ), .S(n8433), .Y(n7758) );
  MUX2X1 U10917 ( .B(\RF[16][46] ), .A(\RF[17][46] ), .S(n8433), .Y(n7757) );
  MUX2X1 U10918 ( .B(n7756), .A(n7753), .S(n8531), .Y(n7760) );
  MUX2X1 U10919 ( .B(\RF[14][46] ), .A(\RF[15][46] ), .S(n8433), .Y(n7764) );
  MUX2X1 U10920 ( .B(\RF[12][46] ), .A(\RF[13][46] ), .S(n8433), .Y(n7763) );
  MUX2X1 U10921 ( .B(\RF[10][46] ), .A(\RF[11][46] ), .S(n8433), .Y(n7767) );
  MUX2X1 U10922 ( .B(\RF[8][46] ), .A(\RF[9][46] ), .S(n8433), .Y(n7766) );
  MUX2X1 U10923 ( .B(n7765), .A(n7762), .S(n8531), .Y(n7776) );
  MUX2X1 U10924 ( .B(\RF[6][46] ), .A(\RF[7][46] ), .S(n8434), .Y(n7770) );
  MUX2X1 U10925 ( .B(\RF[4][46] ), .A(\RF[5][46] ), .S(n8434), .Y(n7769) );
  MUX2X1 U10926 ( .B(\RF[2][46] ), .A(\RF[3][46] ), .S(n8434), .Y(n7773) );
  MUX2X1 U10927 ( .B(\RF[0][46] ), .A(\RF[1][46] ), .S(n8434), .Y(n7772) );
  MUX2X1 U10928 ( .B(n7771), .A(n7768), .S(n8531), .Y(n7775) );
  MUX2X1 U10929 ( .B(n7774), .A(n7759), .S(N17), .Y(n8333) );
  MUX2X1 U10930 ( .B(\RF[30][47] ), .A(\RF[31][47] ), .S(n8434), .Y(n7779) );
  MUX2X1 U10931 ( .B(\RF[28][47] ), .A(\RF[29][47] ), .S(n8434), .Y(n7778) );
  MUX2X1 U10932 ( .B(\RF[26][47] ), .A(\RF[27][47] ), .S(n8434), .Y(n7782) );
  MUX2X1 U10933 ( .B(\RF[24][47] ), .A(\RF[25][47] ), .S(n8434), .Y(n7781) );
  MUX2X1 U10934 ( .B(n7780), .A(n7777), .S(n8531), .Y(n7791) );
  MUX2X1 U10935 ( .B(\RF[22][47] ), .A(\RF[23][47] ), .S(n8434), .Y(n7785) );
  MUX2X1 U10936 ( .B(\RF[20][47] ), .A(\RF[21][47] ), .S(n8434), .Y(n7784) );
  MUX2X1 U10937 ( .B(\RF[18][47] ), .A(\RF[19][47] ), .S(n8434), .Y(n7788) );
  MUX2X1 U10938 ( .B(\RF[16][47] ), .A(\RF[17][47] ), .S(n8434), .Y(n7787) );
  MUX2X1 U10939 ( .B(n7786), .A(n7783), .S(n8531), .Y(n7790) );
  MUX2X1 U10940 ( .B(\RF[14][47] ), .A(\RF[15][47] ), .S(n8435), .Y(n7794) );
  MUX2X1 U10941 ( .B(\RF[12][47] ), .A(\RF[13][47] ), .S(n8435), .Y(n7793) );
  MUX2X1 U10942 ( .B(\RF[10][47] ), .A(\RF[11][47] ), .S(n8435), .Y(n7797) );
  MUX2X1 U10943 ( .B(\RF[8][47] ), .A(\RF[9][47] ), .S(n8435), .Y(n7796) );
  MUX2X1 U10944 ( .B(n7795), .A(n7792), .S(n8531), .Y(n7806) );
  MUX2X1 U10945 ( .B(\RF[6][47] ), .A(\RF[7][47] ), .S(n8435), .Y(n7800) );
  MUX2X1 U10946 ( .B(\RF[4][47] ), .A(\RF[5][47] ), .S(n8435), .Y(n7799) );
  MUX2X1 U10947 ( .B(\RF[2][47] ), .A(\RF[3][47] ), .S(n8435), .Y(n7803) );
  MUX2X1 U10948 ( .B(\RF[0][47] ), .A(\RF[1][47] ), .S(n8435), .Y(n7802) );
  MUX2X1 U10949 ( .B(n7801), .A(n7798), .S(n8531), .Y(n7805) );
  MUX2X1 U10950 ( .B(n7804), .A(n7789), .S(N17), .Y(n8334) );
  MUX2X1 U10951 ( .B(\RF[30][48] ), .A(\RF[31][48] ), .S(n8435), .Y(n7809) );
  MUX2X1 U10952 ( .B(\RF[28][48] ), .A(\RF[29][48] ), .S(n8435), .Y(n7808) );
  MUX2X1 U10953 ( .B(\RF[26][48] ), .A(\RF[27][48] ), .S(n8435), .Y(n7812) );
  MUX2X1 U10954 ( .B(\RF[24][48] ), .A(\RF[25][48] ), .S(n8435), .Y(n7811) );
  MUX2X1 U10955 ( .B(n7810), .A(n7807), .S(n8531), .Y(n7821) );
  MUX2X1 U10956 ( .B(\RF[22][48] ), .A(\RF[23][48] ), .S(n8436), .Y(n7815) );
  MUX2X1 U10957 ( .B(\RF[20][48] ), .A(\RF[21][48] ), .S(n8436), .Y(n7814) );
  MUX2X1 U10958 ( .B(\RF[18][48] ), .A(\RF[19][48] ), .S(n8436), .Y(n7818) );
  MUX2X1 U10959 ( .B(\RF[16][48] ), .A(\RF[17][48] ), .S(n8436), .Y(n7817) );
  MUX2X1 U10960 ( .B(n7816), .A(n7813), .S(n8531), .Y(n7820) );
  MUX2X1 U10961 ( .B(\RF[14][48] ), .A(\RF[15][48] ), .S(n8436), .Y(n7824) );
  MUX2X1 U10962 ( .B(\RF[12][48] ), .A(\RF[13][48] ), .S(n8436), .Y(n7823) );
  MUX2X1 U10963 ( .B(\RF[10][48] ), .A(\RF[11][48] ), .S(n8436), .Y(n7827) );
  MUX2X1 U10964 ( .B(\RF[8][48] ), .A(\RF[9][48] ), .S(n8436), .Y(n7826) );
  MUX2X1 U10965 ( .B(n7825), .A(n7822), .S(n8531), .Y(n7836) );
  MUX2X1 U10966 ( .B(\RF[6][48] ), .A(\RF[7][48] ), .S(n8436), .Y(n7830) );
  MUX2X1 U10967 ( .B(\RF[4][48] ), .A(\RF[5][48] ), .S(n8436), .Y(n7829) );
  MUX2X1 U10968 ( .B(\RF[2][48] ), .A(\RF[3][48] ), .S(n8436), .Y(n7833) );
  MUX2X1 U10969 ( .B(\RF[0][48] ), .A(\RF[1][48] ), .S(n8436), .Y(n7832) );
  MUX2X1 U10970 ( .B(n7831), .A(n7828), .S(n8531), .Y(n7835) );
  MUX2X1 U10971 ( .B(n7834), .A(n7819), .S(N17), .Y(n8335) );
  MUX2X1 U10972 ( .B(\RF[30][49] ), .A(\RF[31][49] ), .S(n8437), .Y(n7839) );
  MUX2X1 U10973 ( .B(\RF[28][49] ), .A(\RF[29][49] ), .S(n8437), .Y(n7838) );
  MUX2X1 U10974 ( .B(\RF[26][49] ), .A(\RF[27][49] ), .S(n8437), .Y(n7842) );
  MUX2X1 U10975 ( .B(\RF[24][49] ), .A(\RF[25][49] ), .S(n8437), .Y(n7841) );
  MUX2X1 U10976 ( .B(n7840), .A(n7837), .S(n8527), .Y(n7851) );
  MUX2X1 U10977 ( .B(\RF[22][49] ), .A(\RF[23][49] ), .S(n8437), .Y(n7845) );
  MUX2X1 U10978 ( .B(\RF[20][49] ), .A(\RF[21][49] ), .S(n8437), .Y(n7844) );
  MUX2X1 U10979 ( .B(\RF[18][49] ), .A(\RF[19][49] ), .S(n8437), .Y(n7848) );
  MUX2X1 U10980 ( .B(\RF[16][49] ), .A(\RF[17][49] ), .S(n8437), .Y(n7847) );
  MUX2X1 U10981 ( .B(n7846), .A(n7843), .S(n8521), .Y(n7850) );
  MUX2X1 U10982 ( .B(\RF[14][49] ), .A(\RF[15][49] ), .S(n8437), .Y(n7854) );
  MUX2X1 U10983 ( .B(\RF[12][49] ), .A(\RF[13][49] ), .S(n8437), .Y(n7853) );
  MUX2X1 U10984 ( .B(\RF[10][49] ), .A(\RF[11][49] ), .S(n8437), .Y(n7857) );
  MUX2X1 U10985 ( .B(\RF[8][49] ), .A(\RF[9][49] ), .S(n8437), .Y(n7856) );
  MUX2X1 U10986 ( .B(n7855), .A(n7852), .S(n8523), .Y(n7866) );
  MUX2X1 U10987 ( .B(\RF[6][49] ), .A(\RF[7][49] ), .S(n8438), .Y(n7860) );
  MUX2X1 U10988 ( .B(\RF[4][49] ), .A(\RF[5][49] ), .S(n8438), .Y(n7859) );
  MUX2X1 U10989 ( .B(\RF[2][49] ), .A(\RF[3][49] ), .S(n8438), .Y(n7863) );
  MUX2X1 U10990 ( .B(\RF[0][49] ), .A(\RF[1][49] ), .S(n8438), .Y(n7862) );
  MUX2X1 U10991 ( .B(n7861), .A(n7858), .S(n8524), .Y(n7865) );
  MUX2X1 U10992 ( .B(n7864), .A(n7849), .S(N17), .Y(n8336) );
  MUX2X1 U10993 ( .B(\RF[30][50] ), .A(\RF[31][50] ), .S(n8438), .Y(n7869) );
  MUX2X1 U10994 ( .B(\RF[28][50] ), .A(\RF[29][50] ), .S(n8438), .Y(n7868) );
  MUX2X1 U10995 ( .B(\RF[26][50] ), .A(\RF[27][50] ), .S(n8438), .Y(n7872) );
  MUX2X1 U10996 ( .B(\RF[24][50] ), .A(\RF[25][50] ), .S(n8438), .Y(n7871) );
  MUX2X1 U10997 ( .B(n7870), .A(n7867), .S(n8529), .Y(n7881) );
  MUX2X1 U10998 ( .B(\RF[22][50] ), .A(\RF[23][50] ), .S(n8438), .Y(n7875) );
  MUX2X1 U10999 ( .B(\RF[20][50] ), .A(\RF[21][50] ), .S(n8438), .Y(n7874) );
  MUX2X1 U11000 ( .B(\RF[18][50] ), .A(\RF[19][50] ), .S(n8438), .Y(n7878) );
  MUX2X1 U11001 ( .B(\RF[16][50] ), .A(\RF[17][50] ), .S(n8438), .Y(n7877) );
  MUX2X1 U11002 ( .B(n7876), .A(n7873), .S(n8519), .Y(n7880) );
  MUX2X1 U11003 ( .B(\RF[14][50] ), .A(\RF[15][50] ), .S(n8439), .Y(n7884) );
  MUX2X1 U11004 ( .B(\RF[12][50] ), .A(\RF[13][50] ), .S(n8439), .Y(n7883) );
  MUX2X1 U11005 ( .B(\RF[10][50] ), .A(\RF[11][50] ), .S(n8439), .Y(n7887) );
  MUX2X1 U11006 ( .B(\RF[8][50] ), .A(\RF[9][50] ), .S(n8439), .Y(n7886) );
  MUX2X1 U11007 ( .B(n7885), .A(n7882), .S(n8520), .Y(n7896) );
  MUX2X1 U11008 ( .B(\RF[6][50] ), .A(\RF[7][50] ), .S(n8439), .Y(n7890) );
  MUX2X1 U11009 ( .B(\RF[4][50] ), .A(\RF[5][50] ), .S(n8439), .Y(n7889) );
  MUX2X1 U11010 ( .B(\RF[2][50] ), .A(\RF[3][50] ), .S(n8439), .Y(n7893) );
  MUX2X1 U11011 ( .B(\RF[0][50] ), .A(\RF[1][50] ), .S(n8439), .Y(n7892) );
  MUX2X1 U11012 ( .B(n7891), .A(n7888), .S(N15), .Y(n7895) );
  MUX2X1 U11013 ( .B(n7894), .A(n7879), .S(N17), .Y(n8337) );
  MUX2X1 U11014 ( .B(\RF[30][51] ), .A(\RF[31][51] ), .S(n8439), .Y(n7899) );
  MUX2X1 U11015 ( .B(\RF[28][51] ), .A(\RF[29][51] ), .S(n8439), .Y(n7898) );
  MUX2X1 U11016 ( .B(\RF[26][51] ), .A(\RF[27][51] ), .S(n8439), .Y(n7902) );
  MUX2X1 U11017 ( .B(\RF[24][51] ), .A(\RF[25][51] ), .S(n8439), .Y(n7901) );
  MUX2X1 U11018 ( .B(n7900), .A(n7897), .S(n8525), .Y(n7911) );
  MUX2X1 U11019 ( .B(\RF[22][51] ), .A(\RF[23][51] ), .S(n8440), .Y(n7905) );
  MUX2X1 U11020 ( .B(\RF[20][51] ), .A(\RF[21][51] ), .S(n8440), .Y(n7904) );
  MUX2X1 U11021 ( .B(\RF[18][51] ), .A(\RF[19][51] ), .S(n8440), .Y(n7908) );
  MUX2X1 U11022 ( .B(\RF[16][51] ), .A(\RF[17][51] ), .S(n8440), .Y(n7907) );
  MUX2X1 U11023 ( .B(n7906), .A(n7903), .S(n8530), .Y(n7910) );
  MUX2X1 U11024 ( .B(\RF[14][51] ), .A(\RF[15][51] ), .S(n8440), .Y(n7914) );
  MUX2X1 U11025 ( .B(\RF[12][51] ), .A(\RF[13][51] ), .S(n8440), .Y(n7913) );
  MUX2X1 U11026 ( .B(\RF[10][51] ), .A(\RF[11][51] ), .S(n8440), .Y(n7917) );
  MUX2X1 U11027 ( .B(\RF[8][51] ), .A(\RF[9][51] ), .S(n8440), .Y(n7916) );
  MUX2X1 U11028 ( .B(n7915), .A(n7912), .S(n8522), .Y(n7926) );
  MUX2X1 U11029 ( .B(\RF[6][51] ), .A(\RF[7][51] ), .S(n8440), .Y(n7920) );
  MUX2X1 U11030 ( .B(\RF[4][51] ), .A(\RF[5][51] ), .S(n8440), .Y(n7919) );
  MUX2X1 U11031 ( .B(\RF[2][51] ), .A(\RF[3][51] ), .S(n8440), .Y(n7923) );
  MUX2X1 U11032 ( .B(\RF[0][51] ), .A(\RF[1][51] ), .S(n8440), .Y(n7922) );
  MUX2X1 U11033 ( .B(n7921), .A(n7918), .S(n8531), .Y(n7925) );
  MUX2X1 U11034 ( .B(n7924), .A(n7909), .S(N17), .Y(n8338) );
  MUX2X1 U11035 ( .B(\RF[30][52] ), .A(\RF[31][52] ), .S(n8441), .Y(n7929) );
  MUX2X1 U11036 ( .B(\RF[28][52] ), .A(\RF[29][52] ), .S(n8441), .Y(n7928) );
  MUX2X1 U11037 ( .B(\RF[26][52] ), .A(\RF[27][52] ), .S(n8441), .Y(n7932) );
  MUX2X1 U11038 ( .B(\RF[24][52] ), .A(\RF[25][52] ), .S(n8441), .Y(n7931) );
  MUX2X1 U11039 ( .B(n7930), .A(n7927), .S(n8532), .Y(n7941) );
  MUX2X1 U11040 ( .B(\RF[22][52] ), .A(\RF[23][52] ), .S(n8441), .Y(n7935) );
  MUX2X1 U11041 ( .B(\RF[20][52] ), .A(\RF[21][52] ), .S(n8441), .Y(n7934) );
  MUX2X1 U11042 ( .B(\RF[18][52] ), .A(\RF[19][52] ), .S(n8441), .Y(n7938) );
  MUX2X1 U11043 ( .B(\RF[16][52] ), .A(\RF[17][52] ), .S(n8441), .Y(n7937) );
  MUX2X1 U11044 ( .B(n7936), .A(n7933), .S(n8532), .Y(n7940) );
  MUX2X1 U11045 ( .B(\RF[14][52] ), .A(\RF[15][52] ), .S(n8441), .Y(n7944) );
  MUX2X1 U11046 ( .B(\RF[12][52] ), .A(\RF[13][52] ), .S(n8441), .Y(n7943) );
  MUX2X1 U11047 ( .B(\RF[10][52] ), .A(\RF[11][52] ), .S(n8441), .Y(n7947) );
  MUX2X1 U11048 ( .B(\RF[8][52] ), .A(\RF[9][52] ), .S(n8441), .Y(n7946) );
  MUX2X1 U11049 ( .B(n7945), .A(n7942), .S(n8532), .Y(n7956) );
  MUX2X1 U11050 ( .B(\RF[6][52] ), .A(\RF[7][52] ), .S(n8442), .Y(n7950) );
  MUX2X1 U11051 ( .B(\RF[4][52] ), .A(\RF[5][52] ), .S(n8442), .Y(n7949) );
  MUX2X1 U11052 ( .B(\RF[2][52] ), .A(\RF[3][52] ), .S(n8442), .Y(n7953) );
  MUX2X1 U11053 ( .B(\RF[0][52] ), .A(\RF[1][52] ), .S(n8442), .Y(n7952) );
  MUX2X1 U11054 ( .B(n7951), .A(n7948), .S(n8532), .Y(n7955) );
  MUX2X1 U11055 ( .B(n7954), .A(n7939), .S(N17), .Y(n8339) );
  MUX2X1 U11056 ( .B(\RF[30][53] ), .A(\RF[31][53] ), .S(n8442), .Y(n7959) );
  MUX2X1 U11057 ( .B(\RF[28][53] ), .A(\RF[29][53] ), .S(n8442), .Y(n7958) );
  MUX2X1 U11058 ( .B(\RF[26][53] ), .A(\RF[27][53] ), .S(n8442), .Y(n7962) );
  MUX2X1 U11059 ( .B(\RF[24][53] ), .A(\RF[25][53] ), .S(n8442), .Y(n7961) );
  MUX2X1 U11060 ( .B(n7960), .A(n7957), .S(n8532), .Y(n7971) );
  MUX2X1 U11061 ( .B(\RF[22][53] ), .A(\RF[23][53] ), .S(n8442), .Y(n7965) );
  MUX2X1 U11062 ( .B(\RF[20][53] ), .A(\RF[21][53] ), .S(n8442), .Y(n7964) );
  MUX2X1 U11063 ( .B(\RF[18][53] ), .A(\RF[19][53] ), .S(n8442), .Y(n7968) );
  MUX2X1 U11064 ( .B(\RF[16][53] ), .A(\RF[17][53] ), .S(n8442), .Y(n7967) );
  MUX2X1 U11065 ( .B(n7966), .A(n7963), .S(n8532), .Y(n7970) );
  MUX2X1 U11066 ( .B(\RF[14][53] ), .A(\RF[15][53] ), .S(n8443), .Y(n7974) );
  MUX2X1 U11067 ( .B(\RF[12][53] ), .A(\RF[13][53] ), .S(n8443), .Y(n7973) );
  MUX2X1 U11068 ( .B(\RF[10][53] ), .A(\RF[11][53] ), .S(n8443), .Y(n7977) );
  MUX2X1 U11069 ( .B(\RF[8][53] ), .A(\RF[9][53] ), .S(n8443), .Y(n7976) );
  MUX2X1 U11070 ( .B(n7975), .A(n7972), .S(n8532), .Y(n7986) );
  MUX2X1 U11071 ( .B(\RF[6][53] ), .A(\RF[7][53] ), .S(n8443), .Y(n7980) );
  MUX2X1 U11072 ( .B(\RF[4][53] ), .A(\RF[5][53] ), .S(n8443), .Y(n7979) );
  MUX2X1 U11073 ( .B(\RF[2][53] ), .A(\RF[3][53] ), .S(n8443), .Y(n7983) );
  MUX2X1 U11074 ( .B(\RF[0][53] ), .A(\RF[1][53] ), .S(n8443), .Y(n7982) );
  MUX2X1 U11075 ( .B(n7981), .A(n7978), .S(n8532), .Y(n7985) );
  MUX2X1 U11076 ( .B(n7984), .A(n7969), .S(N17), .Y(n8340) );
  MUX2X1 U11077 ( .B(\RF[30][54] ), .A(\RF[31][54] ), .S(n8443), .Y(n7989) );
  MUX2X1 U11078 ( .B(\RF[28][54] ), .A(\RF[29][54] ), .S(n8443), .Y(n7988) );
  MUX2X1 U11079 ( .B(\RF[26][54] ), .A(\RF[27][54] ), .S(n8443), .Y(n7992) );
  MUX2X1 U11080 ( .B(\RF[24][54] ), .A(\RF[25][54] ), .S(n8443), .Y(n7991) );
  MUX2X1 U11081 ( .B(n7990), .A(n7987), .S(n8532), .Y(n8001) );
  MUX2X1 U11082 ( .B(\RF[22][54] ), .A(\RF[23][54] ), .S(n8444), .Y(n7995) );
  MUX2X1 U11083 ( .B(\RF[20][54] ), .A(\RF[21][54] ), .S(n8444), .Y(n7994) );
  MUX2X1 U11084 ( .B(\RF[18][54] ), .A(\RF[19][54] ), .S(n8444), .Y(n7998) );
  MUX2X1 U11085 ( .B(\RF[16][54] ), .A(\RF[17][54] ), .S(n8444), .Y(n7997) );
  MUX2X1 U11086 ( .B(n7996), .A(n7993), .S(n8532), .Y(n8000) );
  MUX2X1 U11087 ( .B(\RF[14][54] ), .A(\RF[15][54] ), .S(n8444), .Y(n8004) );
  MUX2X1 U11088 ( .B(\RF[12][54] ), .A(\RF[13][54] ), .S(n8444), .Y(n8003) );
  MUX2X1 U11089 ( .B(\RF[10][54] ), .A(\RF[11][54] ), .S(n8444), .Y(n8007) );
  MUX2X1 U11090 ( .B(\RF[8][54] ), .A(\RF[9][54] ), .S(n8444), .Y(n8006) );
  MUX2X1 U11091 ( .B(n8005), .A(n8002), .S(n8532), .Y(n8016) );
  MUX2X1 U11092 ( .B(\RF[6][54] ), .A(\RF[7][54] ), .S(n8444), .Y(n8010) );
  MUX2X1 U11093 ( .B(\RF[4][54] ), .A(\RF[5][54] ), .S(n8444), .Y(n8009) );
  MUX2X1 U11094 ( .B(\RF[2][54] ), .A(\RF[3][54] ), .S(n8444), .Y(n8013) );
  MUX2X1 U11095 ( .B(\RF[0][54] ), .A(\RF[1][54] ), .S(n8444), .Y(n8012) );
  MUX2X1 U11096 ( .B(n8011), .A(n8008), .S(n8532), .Y(n8015) );
  MUX2X1 U11097 ( .B(n8014), .A(n7999), .S(N17), .Y(n8341) );
  MUX2X1 U11098 ( .B(\RF[30][55] ), .A(\RF[31][55] ), .S(n8445), .Y(n8019) );
  MUX2X1 U11099 ( .B(\RF[28][55] ), .A(\RF[29][55] ), .S(n8445), .Y(n8018) );
  MUX2X1 U11100 ( .B(\RF[26][55] ), .A(\RF[27][55] ), .S(n8445), .Y(n8022) );
  MUX2X1 U11101 ( .B(\RF[24][55] ), .A(\RF[25][55] ), .S(n8445), .Y(n8021) );
  MUX2X1 U11102 ( .B(n8020), .A(n8017), .S(n8533), .Y(n8031) );
  MUX2X1 U11103 ( .B(\RF[22][55] ), .A(\RF[23][55] ), .S(n8445), .Y(n8025) );
  MUX2X1 U11104 ( .B(\RF[20][55] ), .A(\RF[21][55] ), .S(n8445), .Y(n8024) );
  MUX2X1 U11105 ( .B(\RF[18][55] ), .A(\RF[19][55] ), .S(n8445), .Y(n8028) );
  MUX2X1 U11106 ( .B(\RF[16][55] ), .A(\RF[17][55] ), .S(n8445), .Y(n8027) );
  MUX2X1 U11107 ( .B(n8026), .A(n8023), .S(n8533), .Y(n8030) );
  MUX2X1 U11108 ( .B(\RF[14][55] ), .A(\RF[15][55] ), .S(n8445), .Y(n8034) );
  MUX2X1 U11109 ( .B(\RF[12][55] ), .A(\RF[13][55] ), .S(n8445), .Y(n8033) );
  MUX2X1 U11110 ( .B(\RF[10][55] ), .A(\RF[11][55] ), .S(n8445), .Y(n8037) );
  MUX2X1 U11111 ( .B(\RF[8][55] ), .A(\RF[9][55] ), .S(n8445), .Y(n8036) );
  MUX2X1 U11112 ( .B(n8035), .A(n8032), .S(n8533), .Y(n8046) );
  MUX2X1 U11113 ( .B(\RF[6][55] ), .A(\RF[7][55] ), .S(n8446), .Y(n8040) );
  MUX2X1 U11114 ( .B(\RF[4][55] ), .A(\RF[5][55] ), .S(n8446), .Y(n8039) );
  MUX2X1 U11115 ( .B(\RF[2][55] ), .A(\RF[3][55] ), .S(n8446), .Y(n8043) );
  MUX2X1 U11116 ( .B(\RF[0][55] ), .A(\RF[1][55] ), .S(n8446), .Y(n8042) );
  MUX2X1 U11117 ( .B(n8041), .A(n8038), .S(n8533), .Y(n8045) );
  MUX2X1 U11118 ( .B(n8044), .A(n8029), .S(N17), .Y(n8342) );
  MUX2X1 U11119 ( .B(\RF[30][56] ), .A(\RF[31][56] ), .S(n8446), .Y(n8049) );
  MUX2X1 U11120 ( .B(\RF[28][56] ), .A(\RF[29][56] ), .S(n8446), .Y(n8048) );
  MUX2X1 U11121 ( .B(\RF[26][56] ), .A(\RF[27][56] ), .S(n8446), .Y(n8052) );
  MUX2X1 U11122 ( .B(\RF[24][56] ), .A(\RF[25][56] ), .S(n8446), .Y(n8051) );
  MUX2X1 U11123 ( .B(n8050), .A(n8047), .S(n8533), .Y(n8061) );
  MUX2X1 U11124 ( .B(\RF[22][56] ), .A(\RF[23][56] ), .S(n8446), .Y(n8055) );
  MUX2X1 U11125 ( .B(\RF[20][56] ), .A(\RF[21][56] ), .S(n8446), .Y(n8054) );
  MUX2X1 U11126 ( .B(\RF[18][56] ), .A(\RF[19][56] ), .S(n8446), .Y(n8058) );
  MUX2X1 U11127 ( .B(\RF[16][56] ), .A(\RF[17][56] ), .S(n8446), .Y(n8057) );
  MUX2X1 U11128 ( .B(n8056), .A(n8053), .S(n8533), .Y(n8060) );
  MUX2X1 U11129 ( .B(\RF[14][56] ), .A(\RF[15][56] ), .S(n8447), .Y(n8064) );
  MUX2X1 U11130 ( .B(\RF[12][56] ), .A(\RF[13][56] ), .S(n8447), .Y(n8063) );
  MUX2X1 U11131 ( .B(\RF[10][56] ), .A(\RF[11][56] ), .S(n8447), .Y(n8067) );
  MUX2X1 U11132 ( .B(\RF[8][56] ), .A(\RF[9][56] ), .S(n8447), .Y(n8066) );
  MUX2X1 U11133 ( .B(n8065), .A(n8062), .S(n8533), .Y(n8076) );
  MUX2X1 U11134 ( .B(\RF[6][56] ), .A(\RF[7][56] ), .S(n8447), .Y(n8070) );
  MUX2X1 U11135 ( .B(\RF[4][56] ), .A(\RF[5][56] ), .S(n8447), .Y(n8069) );
  MUX2X1 U11136 ( .B(\RF[2][56] ), .A(\RF[3][56] ), .S(n8447), .Y(n8073) );
  MUX2X1 U11137 ( .B(\RF[0][56] ), .A(\RF[1][56] ), .S(n8447), .Y(n8072) );
  MUX2X1 U11138 ( .B(n8071), .A(n8068), .S(n8533), .Y(n8075) );
  MUX2X1 U11139 ( .B(n8074), .A(n8059), .S(N17), .Y(n8343) );
  MUX2X1 U11140 ( .B(\RF[30][57] ), .A(\RF[31][57] ), .S(n8447), .Y(n8079) );
  MUX2X1 U11141 ( .B(\RF[28][57] ), .A(\RF[29][57] ), .S(n8447), .Y(n8078) );
  MUX2X1 U11142 ( .B(\RF[26][57] ), .A(\RF[27][57] ), .S(n8447), .Y(n8082) );
  MUX2X1 U11143 ( .B(\RF[24][57] ), .A(\RF[25][57] ), .S(n8447), .Y(n8081) );
  MUX2X1 U11144 ( .B(n8080), .A(n8077), .S(n8533), .Y(n8091) );
  MUX2X1 U11145 ( .B(\RF[22][57] ), .A(\RF[23][57] ), .S(n8448), .Y(n8085) );
  MUX2X1 U11146 ( .B(\RF[20][57] ), .A(\RF[21][57] ), .S(n8448), .Y(n8084) );
  MUX2X1 U11147 ( .B(\RF[18][57] ), .A(\RF[19][57] ), .S(n8448), .Y(n8088) );
  MUX2X1 U11148 ( .B(\RF[16][57] ), .A(\RF[17][57] ), .S(n8448), .Y(n8087) );
  MUX2X1 U11149 ( .B(n8086), .A(n8083), .S(n8533), .Y(n8090) );
  MUX2X1 U11150 ( .B(\RF[14][57] ), .A(\RF[15][57] ), .S(n8448), .Y(n8094) );
  MUX2X1 U11151 ( .B(\RF[12][57] ), .A(\RF[13][57] ), .S(n8448), .Y(n8093) );
  MUX2X1 U11152 ( .B(\RF[10][57] ), .A(\RF[11][57] ), .S(n8448), .Y(n8097) );
  MUX2X1 U11153 ( .B(\RF[8][57] ), .A(\RF[9][57] ), .S(n8448), .Y(n8096) );
  MUX2X1 U11154 ( .B(n8095), .A(n8092), .S(n8533), .Y(n8106) );
  MUX2X1 U11155 ( .B(\RF[6][57] ), .A(\RF[7][57] ), .S(n8448), .Y(n8100) );
  MUX2X1 U11156 ( .B(\RF[4][57] ), .A(\RF[5][57] ), .S(n8448), .Y(n8099) );
  MUX2X1 U11157 ( .B(\RF[2][57] ), .A(\RF[3][57] ), .S(n8448), .Y(n8103) );
  MUX2X1 U11158 ( .B(\RF[0][57] ), .A(\RF[1][57] ), .S(n8448), .Y(n8102) );
  MUX2X1 U11159 ( .B(n8101), .A(n8098), .S(n8533), .Y(n8105) );
  MUX2X1 U11160 ( .B(n8104), .A(n8089), .S(N17), .Y(n8344) );
  MUX2X1 U11161 ( .B(\RF[30][58] ), .A(\RF[31][58] ), .S(n8449), .Y(n8109) );
  MUX2X1 U11162 ( .B(\RF[28][58] ), .A(\RF[29][58] ), .S(n8449), .Y(n8108) );
  MUX2X1 U11163 ( .B(\RF[26][58] ), .A(\RF[27][58] ), .S(n8449), .Y(n8112) );
  MUX2X1 U11164 ( .B(\RF[24][58] ), .A(\RF[25][58] ), .S(n8449), .Y(n8111) );
  MUX2X1 U11165 ( .B(n8110), .A(n8107), .S(n8526), .Y(n8121) );
  MUX2X1 U11166 ( .B(\RF[22][58] ), .A(\RF[23][58] ), .S(n8449), .Y(n8115) );
  MUX2X1 U11167 ( .B(\RF[20][58] ), .A(\RF[21][58] ), .S(n8449), .Y(n8114) );
  MUX2X1 U11168 ( .B(\RF[18][58] ), .A(\RF[19][58] ), .S(n8449), .Y(n8118) );
  MUX2X1 U11169 ( .B(\RF[16][58] ), .A(\RF[17][58] ), .S(n8449), .Y(n8117) );
  MUX2X1 U11170 ( .B(n8116), .A(n8113), .S(n8528), .Y(n8120) );
  MUX2X1 U11171 ( .B(\RF[14][58] ), .A(\RF[15][58] ), .S(n8449), .Y(n8124) );
  MUX2X1 U11172 ( .B(\RF[12][58] ), .A(\RF[13][58] ), .S(n8449), .Y(n8123) );
  MUX2X1 U11173 ( .B(\RF[10][58] ), .A(\RF[11][58] ), .S(n8449), .Y(n8127) );
  MUX2X1 U11174 ( .B(\RF[8][58] ), .A(\RF[9][58] ), .S(n8449), .Y(n8126) );
  MUX2X1 U11175 ( .B(n8125), .A(n8122), .S(n8532), .Y(n8136) );
  MUX2X1 U11176 ( .B(\RF[6][58] ), .A(\RF[7][58] ), .S(n8450), .Y(n8130) );
  MUX2X1 U11177 ( .B(\RF[4][58] ), .A(\RF[5][58] ), .S(n8450), .Y(n8129) );
  MUX2X1 U11178 ( .B(\RF[2][58] ), .A(\RF[3][58] ), .S(n8450), .Y(n8133) );
  MUX2X1 U11179 ( .B(\RF[0][58] ), .A(\RF[1][58] ), .S(n8450), .Y(n8132) );
  MUX2X1 U11180 ( .B(n8131), .A(n8128), .S(n8533), .Y(n8135) );
  MUX2X1 U11181 ( .B(n8134), .A(n8119), .S(N17), .Y(n8345) );
  MUX2X1 U11182 ( .B(\RF[30][59] ), .A(\RF[31][59] ), .S(n8450), .Y(n8139) );
  MUX2X1 U11183 ( .B(\RF[28][59] ), .A(\RF[29][59] ), .S(n8450), .Y(n8138) );
  MUX2X1 U11184 ( .B(\RF[26][59] ), .A(\RF[27][59] ), .S(n8450), .Y(n8142) );
  MUX2X1 U11185 ( .B(\RF[24][59] ), .A(\RF[25][59] ), .S(n8450), .Y(n8141) );
  MUX2X1 U11186 ( .B(n8140), .A(n8137), .S(n8517), .Y(n8151) );
  MUX2X1 U11187 ( .B(\RF[22][59] ), .A(\RF[23][59] ), .S(n8450), .Y(n8145) );
  MUX2X1 U11188 ( .B(\RF[20][59] ), .A(\RF[21][59] ), .S(n8450), .Y(n8144) );
  MUX2X1 U11189 ( .B(\RF[18][59] ), .A(\RF[19][59] ), .S(n8450), .Y(n8148) );
  MUX2X1 U11190 ( .B(\RF[16][59] ), .A(\RF[17][59] ), .S(n8450), .Y(n8147) );
  MUX2X1 U11191 ( .B(n8146), .A(n8143), .S(n8518), .Y(n8150) );
  MUX2X1 U11192 ( .B(\RF[14][59] ), .A(\RF[15][59] ), .S(n8451), .Y(n8154) );
  MUX2X1 U11193 ( .B(\RF[12][59] ), .A(\RF[13][59] ), .S(n8451), .Y(n8153) );
  MUX2X1 U11194 ( .B(\RF[10][59] ), .A(\RF[11][59] ), .S(n8451), .Y(n8157) );
  MUX2X1 U11195 ( .B(\RF[8][59] ), .A(\RF[9][59] ), .S(n8451), .Y(n8156) );
  MUX2X1 U11196 ( .B(n8155), .A(n8152), .S(n8527), .Y(n8166) );
  MUX2X1 U11197 ( .B(\RF[6][59] ), .A(\RF[7][59] ), .S(n8451), .Y(n8160) );
  MUX2X1 U11198 ( .B(\RF[4][59] ), .A(\RF[5][59] ), .S(n8451), .Y(n8159) );
  MUX2X1 U11199 ( .B(\RF[2][59] ), .A(\RF[3][59] ), .S(n8451), .Y(n8163) );
  MUX2X1 U11200 ( .B(\RF[0][59] ), .A(\RF[1][59] ), .S(n8451), .Y(n8162) );
  MUX2X1 U11201 ( .B(n8161), .A(n8158), .S(n8518), .Y(n8165) );
  MUX2X1 U11202 ( .B(n8164), .A(n8149), .S(N17), .Y(n8346) );
  MUX2X1 U11203 ( .B(\RF[30][60] ), .A(\RF[31][60] ), .S(n8451), .Y(n8169) );
  MUX2X1 U11204 ( .B(\RF[28][60] ), .A(\RF[29][60] ), .S(n8451), .Y(n8168) );
  MUX2X1 U11205 ( .B(\RF[26][60] ), .A(\RF[27][60] ), .S(n8451), .Y(n8172) );
  MUX2X1 U11206 ( .B(\RF[24][60] ), .A(\RF[25][60] ), .S(n8451), .Y(n8171) );
  MUX2X1 U11207 ( .B(n8170), .A(n8167), .S(n8521), .Y(n8181) );
  MUX2X1 U11208 ( .B(\RF[22][60] ), .A(\RF[23][60] ), .S(n8452), .Y(n8175) );
  MUX2X1 U11209 ( .B(\RF[20][60] ), .A(\RF[21][60] ), .S(n8452), .Y(n8174) );
  MUX2X1 U11210 ( .B(\RF[18][60] ), .A(\RF[19][60] ), .S(n8452), .Y(n8178) );
  MUX2X1 U11211 ( .B(\RF[16][60] ), .A(\RF[17][60] ), .S(n8452), .Y(n8177) );
  MUX2X1 U11212 ( .B(n8176), .A(n8173), .S(n8523), .Y(n8180) );
  MUX2X1 U11213 ( .B(\RF[14][60] ), .A(\RF[15][60] ), .S(n8452), .Y(n8184) );
  MUX2X1 U11214 ( .B(\RF[12][60] ), .A(\RF[13][60] ), .S(n8452), .Y(n8183) );
  MUX2X1 U11215 ( .B(\RF[10][60] ), .A(\RF[11][60] ), .S(n8452), .Y(n8187) );
  MUX2X1 U11216 ( .B(\RF[8][60] ), .A(\RF[9][60] ), .S(n8452), .Y(n8186) );
  MUX2X1 U11217 ( .B(n8185), .A(n8182), .S(n8524), .Y(n8196) );
  MUX2X1 U11218 ( .B(\RF[6][60] ), .A(\RF[7][60] ), .S(n8452), .Y(n8190) );
  MUX2X1 U11219 ( .B(\RF[4][60] ), .A(\RF[5][60] ), .S(n8452), .Y(n8189) );
  MUX2X1 U11220 ( .B(\RF[2][60] ), .A(\RF[3][60] ), .S(n8452), .Y(n8193) );
  MUX2X1 U11221 ( .B(\RF[0][60] ), .A(\RF[1][60] ), .S(n8452), .Y(n8192) );
  MUX2X1 U11222 ( .B(n8191), .A(n8188), .S(n8529), .Y(n8195) );
  MUX2X1 U11223 ( .B(n8194), .A(n8179), .S(N17), .Y(n8347) );
  MUX2X1 U11224 ( .B(\RF[30][61] ), .A(\RF[31][61] ), .S(n8453), .Y(n8199) );
  MUX2X1 U11225 ( .B(\RF[28][61] ), .A(\RF[29][61] ), .S(n8453), .Y(n8198) );
  MUX2X1 U11226 ( .B(\RF[26][61] ), .A(\RF[27][61] ), .S(n8453), .Y(n8202) );
  MUX2X1 U11227 ( .B(\RF[24][61] ), .A(\RF[25][61] ), .S(n8453), .Y(n8201) );
  MUX2X1 U11228 ( .B(n8200), .A(n8197), .S(N15), .Y(n8211) );
  MUX2X1 U11229 ( .B(\RF[22][61] ), .A(\RF[23][61] ), .S(n8453), .Y(n8205) );
  MUX2X1 U11230 ( .B(\RF[20][61] ), .A(\RF[21][61] ), .S(n8453), .Y(n8204) );
  MUX2X1 U11231 ( .B(\RF[18][61] ), .A(\RF[19][61] ), .S(n8453), .Y(n8208) );
  MUX2X1 U11232 ( .B(\RF[16][61] ), .A(\RF[17][61] ), .S(n8453), .Y(n8207) );
  MUX2X1 U11233 ( .B(n8206), .A(n8203), .S(N15), .Y(n8210) );
  MUX2X1 U11234 ( .B(\RF[14][61] ), .A(\RF[15][61] ), .S(n8453), .Y(n8214) );
  MUX2X1 U11235 ( .B(\RF[12][61] ), .A(\RF[13][61] ), .S(n8453), .Y(n8213) );
  MUX2X1 U11236 ( .B(\RF[10][61] ), .A(\RF[11][61] ), .S(n8453), .Y(n8217) );
  MUX2X1 U11237 ( .B(\RF[8][61] ), .A(\RF[9][61] ), .S(n8453), .Y(n8216) );
  MUX2X1 U11238 ( .B(n8215), .A(n8212), .S(N15), .Y(n8226) );
  MUX2X1 U11239 ( .B(\RF[6][61] ), .A(\RF[7][61] ), .S(n8454), .Y(n8220) );
  MUX2X1 U11240 ( .B(\RF[4][61] ), .A(\RF[5][61] ), .S(n8454), .Y(n8219) );
  MUX2X1 U11241 ( .B(\RF[2][61] ), .A(\RF[3][61] ), .S(n8454), .Y(n8223) );
  MUX2X1 U11242 ( .B(\RF[0][61] ), .A(\RF[1][61] ), .S(n8454), .Y(n8222) );
  MUX2X1 U11243 ( .B(n8221), .A(n8218), .S(N15), .Y(n8225) );
  MUX2X1 U11244 ( .B(n8224), .A(n8209), .S(N17), .Y(n8348) );
  MUX2X1 U11245 ( .B(\RF[30][62] ), .A(\RF[31][62] ), .S(n8454), .Y(n8229) );
  MUX2X1 U11246 ( .B(\RF[28][62] ), .A(\RF[29][62] ), .S(n8454), .Y(n8228) );
  MUX2X1 U11247 ( .B(\RF[26][62] ), .A(\RF[27][62] ), .S(n8454), .Y(n8232) );
  MUX2X1 U11248 ( .B(\RF[24][62] ), .A(\RF[25][62] ), .S(n8454), .Y(n8231) );
  MUX2X1 U11249 ( .B(n8230), .A(n8227), .S(N15), .Y(n8241) );
  MUX2X1 U11250 ( .B(\RF[22][62] ), .A(\RF[23][62] ), .S(n8454), .Y(n8235) );
  MUX2X1 U11251 ( .B(\RF[20][62] ), .A(\RF[21][62] ), .S(n8454), .Y(n8234) );
  MUX2X1 U11252 ( .B(\RF[18][62] ), .A(\RF[19][62] ), .S(n8454), .Y(n8238) );
  MUX2X1 U11253 ( .B(\RF[16][62] ), .A(\RF[17][62] ), .S(n8454), .Y(n8237) );
  MUX2X1 U11254 ( .B(n8236), .A(n8233), .S(N15), .Y(n8240) );
  MUX2X1 U11255 ( .B(\RF[14][62] ), .A(\RF[15][62] ), .S(n8455), .Y(n8244) );
  MUX2X1 U11256 ( .B(\RF[12][62] ), .A(\RF[13][62] ), .S(n8455), .Y(n8243) );
  MUX2X1 U11257 ( .B(\RF[10][62] ), .A(\RF[11][62] ), .S(n8455), .Y(n8247) );
  MUX2X1 U11258 ( .B(\RF[8][62] ), .A(\RF[9][62] ), .S(n8455), .Y(n8246) );
  MUX2X1 U11259 ( .B(n8245), .A(n8242), .S(N15), .Y(n8256) );
  MUX2X1 U11260 ( .B(\RF[6][62] ), .A(\RF[7][62] ), .S(n8455), .Y(n8250) );
  MUX2X1 U11261 ( .B(\RF[4][62] ), .A(\RF[5][62] ), .S(n8455), .Y(n8249) );
  MUX2X1 U11262 ( .B(\RF[2][62] ), .A(\RF[3][62] ), .S(n8455), .Y(n8253) );
  MUX2X1 U11263 ( .B(\RF[0][62] ), .A(\RF[1][62] ), .S(n8455), .Y(n8252) );
  MUX2X1 U11264 ( .B(n8251), .A(n8248), .S(N15), .Y(n8255) );
  MUX2X1 U11265 ( .B(n8254), .A(n8239), .S(N17), .Y(n8349) );
  MUX2X1 U11266 ( .B(\RF[30][63] ), .A(\RF[31][63] ), .S(n8455), .Y(n8259) );
  MUX2X1 U11267 ( .B(\RF[28][63] ), .A(\RF[29][63] ), .S(n8455), .Y(n8258) );
  MUX2X1 U11268 ( .B(\RF[26][63] ), .A(\RF[27][63] ), .S(n8455), .Y(n8262) );
  MUX2X1 U11269 ( .B(\RF[24][63] ), .A(\RF[25][63] ), .S(n8455), .Y(n8261) );
  MUX2X1 U11270 ( .B(n8260), .A(n8257), .S(n8525), .Y(n8271) );
  MUX2X1 U11271 ( .B(\RF[22][63] ), .A(\RF[23][63] ), .S(n8456), .Y(n8265) );
  MUX2X1 U11272 ( .B(\RF[20][63] ), .A(\RF[21][63] ), .S(n8456), .Y(n8264) );
  MUX2X1 U11273 ( .B(\RF[18][63] ), .A(\RF[19][63] ), .S(n8456), .Y(n8268) );
  MUX2X1 U11274 ( .B(\RF[16][63] ), .A(\RF[17][63] ), .S(n8456), .Y(n8267) );
  MUX2X1 U11275 ( .B(n8266), .A(n8263), .S(n8530), .Y(n8270) );
  MUX2X1 U11276 ( .B(\RF[14][63] ), .A(\RF[15][63] ), .S(n8456), .Y(n8274) );
  MUX2X1 U11277 ( .B(\RF[12][63] ), .A(\RF[13][63] ), .S(n8456), .Y(n8273) );
  MUX2X1 U11278 ( .B(\RF[10][63] ), .A(\RF[11][63] ), .S(n8456), .Y(n8277) );
  MUX2X1 U11279 ( .B(\RF[8][63] ), .A(\RF[9][63] ), .S(n8456), .Y(n8276) );
  MUX2X1 U11280 ( .B(n8275), .A(n8272), .S(n8522), .Y(n8286) );
  MUX2X1 U11281 ( .B(\RF[6][63] ), .A(\RF[7][63] ), .S(n8456), .Y(n8280) );
  MUX2X1 U11282 ( .B(\RF[4][63] ), .A(\RF[5][63] ), .S(n8456), .Y(n8279) );
  MUX2X1 U11283 ( .B(\RF[2][63] ), .A(\RF[3][63] ), .S(n8456), .Y(n8283) );
  MUX2X1 U11284 ( .B(\RF[0][63] ), .A(\RF[1][63] ), .S(n8456), .Y(n8282) );
  MUX2X1 U11285 ( .B(n8281), .A(n8278), .S(n8531), .Y(n8285) );
  MUX2X1 U11286 ( .B(n8284), .A(n8269), .S(N17), .Y(n8350) );
  MUX2X1 U11287 ( .B(n8535), .A(n8536), .S(n10639), .Y(n8534) );
  MUX2X1 U11288 ( .B(n8538), .A(n8539), .S(n10639), .Y(n8537) );
  MUX2X1 U11289 ( .B(n8541), .A(n8542), .S(n10639), .Y(n8540) );
  MUX2X1 U11290 ( .B(n8544), .A(n8545), .S(n10639), .Y(n8543) );
  MUX2X1 U11291 ( .B(n8547), .A(n8548), .S(N21), .Y(n8546) );
  MUX2X1 U11292 ( .B(n8550), .A(n8551), .S(n10639), .Y(n8549) );
  MUX2X1 U11293 ( .B(n8553), .A(n8554), .S(n10639), .Y(n8552) );
  MUX2X1 U11294 ( .B(n8556), .A(n8557), .S(n10639), .Y(n8555) );
  MUX2X1 U11295 ( .B(n8559), .A(n8560), .S(n10639), .Y(n8558) );
  MUX2X1 U11296 ( .B(n8562), .A(n8563), .S(N21), .Y(n8561) );
  MUX2X1 U11297 ( .B(n8565), .A(n8566), .S(n10640), .Y(n8564) );
  MUX2X1 U11298 ( .B(n8568), .A(n8569), .S(n10640), .Y(n8567) );
  MUX2X1 U11299 ( .B(n8571), .A(n8572), .S(n10640), .Y(n8570) );
  MUX2X1 U11300 ( .B(n8574), .A(n8575), .S(n10640), .Y(n8573) );
  MUX2X1 U11301 ( .B(n8577), .A(n8578), .S(N21), .Y(n8576) );
  MUX2X1 U11302 ( .B(n8580), .A(n8581), .S(n10640), .Y(n8579) );
  MUX2X1 U11303 ( .B(n8583), .A(n8584), .S(n10640), .Y(n8582) );
  MUX2X1 U11304 ( .B(n8586), .A(n8587), .S(n10640), .Y(n8585) );
  MUX2X1 U11305 ( .B(n8589), .A(n8590), .S(n10640), .Y(n8588) );
  MUX2X1 U11306 ( .B(n8592), .A(n8593), .S(N21), .Y(n8591) );
  MUX2X1 U11307 ( .B(n8595), .A(n8596), .S(n10640), .Y(n8594) );
  MUX2X1 U11308 ( .B(n8598), .A(n8599), .S(n10640), .Y(n8597) );
  MUX2X1 U11309 ( .B(n8601), .A(n8602), .S(n10640), .Y(n8600) );
  MUX2X1 U11310 ( .B(n8604), .A(n8605), .S(n10640), .Y(n8603) );
  MUX2X1 U11311 ( .B(n8607), .A(n8608), .S(N21), .Y(n8606) );
  MUX2X1 U11312 ( .B(n8610), .A(n8611), .S(n10641), .Y(n8609) );
  MUX2X1 U11313 ( .B(n8613), .A(n8614), .S(n10641), .Y(n8612) );
  MUX2X1 U11314 ( .B(n8616), .A(n8617), .S(n10641), .Y(n8615) );
  MUX2X1 U11315 ( .B(n8619), .A(n8620), .S(n10641), .Y(n8618) );
  MUX2X1 U11316 ( .B(n8622), .A(n8623), .S(N21), .Y(n8621) );
  MUX2X1 U11317 ( .B(n8625), .A(n8626), .S(n10641), .Y(n8624) );
  MUX2X1 U11318 ( .B(n8628), .A(n8629), .S(n10641), .Y(n8627) );
  MUX2X1 U11319 ( .B(n8631), .A(n8632), .S(n10641), .Y(n8630) );
  MUX2X1 U11320 ( .B(n8634), .A(n8635), .S(n10641), .Y(n8633) );
  MUX2X1 U11321 ( .B(n8637), .A(n8638), .S(N21), .Y(n8636) );
  MUX2X1 U11322 ( .B(n8640), .A(n8641), .S(n10641), .Y(n8639) );
  MUX2X1 U11323 ( .B(n8643), .A(n8644), .S(n10641), .Y(n8642) );
  MUX2X1 U11324 ( .B(n8646), .A(n8647), .S(n10641), .Y(n8645) );
  MUX2X1 U11325 ( .B(n8649), .A(n8650), .S(n10641), .Y(n8648) );
  MUX2X1 U11326 ( .B(n8652), .A(n8653), .S(N21), .Y(n8651) );
  MUX2X1 U11327 ( .B(n8655), .A(n8656), .S(n10642), .Y(n8654) );
  MUX2X1 U11328 ( .B(n8658), .A(n8659), .S(n10642), .Y(n8657) );
  MUX2X1 U11329 ( .B(n8661), .A(n8662), .S(n10642), .Y(n8660) );
  MUX2X1 U11330 ( .B(n8664), .A(n8665), .S(n10642), .Y(n8663) );
  MUX2X1 U11331 ( .B(n8667), .A(n8668), .S(N21), .Y(n8666) );
  MUX2X1 U11332 ( .B(n8670), .A(n8671), .S(n10642), .Y(n8669) );
  MUX2X1 U11333 ( .B(n8673), .A(n8674), .S(n10642), .Y(n8672) );
  MUX2X1 U11334 ( .B(n8676), .A(n8677), .S(n10642), .Y(n8675) );
  MUX2X1 U11335 ( .B(n8679), .A(n8680), .S(n10642), .Y(n8678) );
  MUX2X1 U11336 ( .B(n8682), .A(n8683), .S(N21), .Y(n8681) );
  MUX2X1 U11337 ( .B(n8685), .A(n8686), .S(n10642), .Y(n8684) );
  MUX2X1 U11338 ( .B(n8688), .A(n8689), .S(n10642), .Y(n8687) );
  MUX2X1 U11339 ( .B(n8691), .A(n8692), .S(n10642), .Y(n8690) );
  MUX2X1 U11340 ( .B(n8694), .A(n8695), .S(n10642), .Y(n8693) );
  MUX2X1 U11341 ( .B(n8697), .A(n8698), .S(N21), .Y(n8696) );
  MUX2X1 U11342 ( .B(n8700), .A(n8701), .S(n10643), .Y(n8699) );
  MUX2X1 U11343 ( .B(n8703), .A(n8704), .S(n10643), .Y(n8702) );
  MUX2X1 U11344 ( .B(n8706), .A(n8707), .S(n10643), .Y(n8705) );
  MUX2X1 U11345 ( .B(n8709), .A(n8710), .S(n10643), .Y(n8708) );
  MUX2X1 U11346 ( .B(n8712), .A(n8713), .S(N21), .Y(n8711) );
  MUX2X1 U11347 ( .B(n8715), .A(n8716), .S(n10643), .Y(n8714) );
  MUX2X1 U11348 ( .B(n8718), .A(n8719), .S(n10643), .Y(n8717) );
  MUX2X1 U11349 ( .B(n8721), .A(n8722), .S(n10643), .Y(n8720) );
  MUX2X1 U11350 ( .B(n8724), .A(n8725), .S(n10643), .Y(n8723) );
  MUX2X1 U11351 ( .B(n8727), .A(n8728), .S(N21), .Y(n8726) );
  MUX2X1 U11352 ( .B(n8730), .A(n8731), .S(n10643), .Y(n8729) );
  MUX2X1 U11353 ( .B(n8733), .A(n8734), .S(n10643), .Y(n8732) );
  MUX2X1 U11354 ( .B(n8736), .A(n8737), .S(n10643), .Y(n8735) );
  MUX2X1 U11355 ( .B(n8739), .A(n8740), .S(n10643), .Y(n8738) );
  MUX2X1 U11356 ( .B(n8742), .A(n8743), .S(N21), .Y(n8741) );
  MUX2X1 U11357 ( .B(n8745), .A(n8746), .S(n10644), .Y(n8744) );
  MUX2X1 U11358 ( .B(n8748), .A(n8749), .S(n10644), .Y(n8747) );
  MUX2X1 U11359 ( .B(n8751), .A(n8752), .S(n10644), .Y(n8750) );
  MUX2X1 U11360 ( .B(n8754), .A(n8755), .S(n10644), .Y(n8753) );
  MUX2X1 U11361 ( .B(n8757), .A(n8758), .S(N21), .Y(n8756) );
  MUX2X1 U11362 ( .B(n8760), .A(n8761), .S(n10644), .Y(n8759) );
  MUX2X1 U11363 ( .B(n8763), .A(n8764), .S(n10644), .Y(n8762) );
  MUX2X1 U11364 ( .B(n8766), .A(n8767), .S(n10644), .Y(n8765) );
  MUX2X1 U11365 ( .B(n8769), .A(n8770), .S(n10644), .Y(n8768) );
  MUX2X1 U11366 ( .B(n8772), .A(n8773), .S(N21), .Y(n8771) );
  MUX2X1 U11367 ( .B(n8775), .A(n8776), .S(n10644), .Y(n8774) );
  MUX2X1 U11368 ( .B(n8778), .A(n8779), .S(n10644), .Y(n8777) );
  MUX2X1 U11369 ( .B(n8781), .A(n8782), .S(n10644), .Y(n8780) );
  MUX2X1 U11370 ( .B(n8784), .A(n8785), .S(n10644), .Y(n8783) );
  MUX2X1 U11371 ( .B(n8787), .A(n8788), .S(N21), .Y(n8786) );
  MUX2X1 U11372 ( .B(n8790), .A(n8791), .S(n10645), .Y(n8789) );
  MUX2X1 U11373 ( .B(n8793), .A(n8794), .S(n10645), .Y(n8792) );
  MUX2X1 U11374 ( .B(n8796), .A(n8797), .S(n10645), .Y(n8795) );
  MUX2X1 U11375 ( .B(n8799), .A(n8800), .S(n10645), .Y(n8798) );
  MUX2X1 U11376 ( .B(n8802), .A(n8803), .S(N21), .Y(n8801) );
  MUX2X1 U11377 ( .B(n8805), .A(n8806), .S(n10645), .Y(n8804) );
  MUX2X1 U11378 ( .B(n8808), .A(n8809), .S(n10645), .Y(n8807) );
  MUX2X1 U11379 ( .B(n8811), .A(n8812), .S(n10645), .Y(n8810) );
  MUX2X1 U11380 ( .B(n8814), .A(n8815), .S(n10645), .Y(n8813) );
  MUX2X1 U11381 ( .B(n8817), .A(n8818), .S(N21), .Y(n8816) );
  MUX2X1 U11382 ( .B(n8820), .A(n8821), .S(n10645), .Y(n8819) );
  MUX2X1 U11383 ( .B(n8823), .A(n8824), .S(n10645), .Y(n8822) );
  MUX2X1 U11384 ( .B(n8826), .A(n8827), .S(n10645), .Y(n8825) );
  MUX2X1 U11385 ( .B(n8829), .A(n8830), .S(n10645), .Y(n8828) );
  MUX2X1 U11386 ( .B(n8832), .A(n8833), .S(N21), .Y(n8831) );
  MUX2X1 U11387 ( .B(n8835), .A(n8836), .S(n10646), .Y(n8834) );
  MUX2X1 U11388 ( .B(n8838), .A(n8839), .S(n10646), .Y(n8837) );
  MUX2X1 U11389 ( .B(n8841), .A(n8842), .S(n10646), .Y(n8840) );
  MUX2X1 U11390 ( .B(n8844), .A(n8845), .S(n10646), .Y(n8843) );
  MUX2X1 U11391 ( .B(n8847), .A(n8848), .S(N21), .Y(n8846) );
  MUX2X1 U11392 ( .B(n8850), .A(n8851), .S(n10646), .Y(n8849) );
  MUX2X1 U11393 ( .B(n8853), .A(n8854), .S(n10646), .Y(n8852) );
  MUX2X1 U11394 ( .B(n8856), .A(n8857), .S(n10646), .Y(n8855) );
  MUX2X1 U11395 ( .B(n8859), .A(n8860), .S(n10646), .Y(n8858) );
  MUX2X1 U11396 ( .B(n8862), .A(n8863), .S(N21), .Y(n8861) );
  MUX2X1 U11397 ( .B(n8865), .A(n8866), .S(n10646), .Y(n8864) );
  MUX2X1 U11398 ( .B(n8868), .A(n8869), .S(n10646), .Y(n8867) );
  MUX2X1 U11399 ( .B(n8871), .A(n8872), .S(n10646), .Y(n8870) );
  MUX2X1 U11400 ( .B(n8874), .A(n8875), .S(n10646), .Y(n8873) );
  MUX2X1 U11401 ( .B(n8877), .A(n8878), .S(N21), .Y(n8876) );
  MUX2X1 U11402 ( .B(n8880), .A(n8881), .S(n10647), .Y(n8879) );
  MUX2X1 U11403 ( .B(n8883), .A(n8884), .S(n10647), .Y(n8882) );
  MUX2X1 U11404 ( .B(n8886), .A(n8887), .S(n10647), .Y(n8885) );
  MUX2X1 U11405 ( .B(n8889), .A(n8890), .S(n10647), .Y(n8888) );
  MUX2X1 U11406 ( .B(n8892), .A(n8893), .S(N21), .Y(n8891) );
  MUX2X1 U11407 ( .B(n8895), .A(n8896), .S(n10647), .Y(n8894) );
  MUX2X1 U11408 ( .B(n8898), .A(n8899), .S(n10647), .Y(n8897) );
  MUX2X1 U11409 ( .B(n8901), .A(n8902), .S(n10647), .Y(n8900) );
  MUX2X1 U11410 ( .B(n8904), .A(n8905), .S(n10647), .Y(n8903) );
  MUX2X1 U11411 ( .B(n8907), .A(n8908), .S(N21), .Y(n8906) );
  MUX2X1 U11412 ( .B(n8910), .A(n8911), .S(n10647), .Y(n8909) );
  MUX2X1 U11413 ( .B(n8913), .A(n8914), .S(n10647), .Y(n8912) );
  MUX2X1 U11414 ( .B(n8916), .A(n8917), .S(n10647), .Y(n8915) );
  MUX2X1 U11415 ( .B(n8919), .A(n8920), .S(n10647), .Y(n8918) );
  MUX2X1 U11416 ( .B(n8922), .A(n8923), .S(N21), .Y(n8921) );
  MUX2X1 U11417 ( .B(n8925), .A(n8926), .S(n10648), .Y(n8924) );
  MUX2X1 U11418 ( .B(n8928), .A(n8929), .S(n10648), .Y(n8927) );
  MUX2X1 U11419 ( .B(n8931), .A(n8932), .S(n10648), .Y(n8930) );
  MUX2X1 U11420 ( .B(n8934), .A(n8935), .S(n10648), .Y(n8933) );
  MUX2X1 U11421 ( .B(n8937), .A(n8938), .S(N21), .Y(n8936) );
  MUX2X1 U11422 ( .B(n8940), .A(n8941), .S(n10648), .Y(n8939) );
  MUX2X1 U11423 ( .B(n8943), .A(n8944), .S(n10648), .Y(n8942) );
  MUX2X1 U11424 ( .B(n8946), .A(n8947), .S(n10648), .Y(n8945) );
  MUX2X1 U11425 ( .B(n8949), .A(n8950), .S(n10648), .Y(n8948) );
  MUX2X1 U11426 ( .B(n8952), .A(n8953), .S(N21), .Y(n8951) );
  MUX2X1 U11427 ( .B(n8955), .A(n8956), .S(n10648), .Y(n8954) );
  MUX2X1 U11428 ( .B(n8958), .A(n8959), .S(n10648), .Y(n8957) );
  MUX2X1 U11429 ( .B(n8961), .A(n8962), .S(n10648), .Y(n8960) );
  MUX2X1 U11430 ( .B(n8964), .A(n8965), .S(n10648), .Y(n8963) );
  MUX2X1 U11431 ( .B(n8967), .A(n8968), .S(N21), .Y(n8966) );
  MUX2X1 U11432 ( .B(n8970), .A(n8971), .S(n10649), .Y(n8969) );
  MUX2X1 U11433 ( .B(n8973), .A(n8974), .S(n10649), .Y(n8972) );
  MUX2X1 U11434 ( .B(n8976), .A(n8977), .S(n10649), .Y(n8975) );
  MUX2X1 U11435 ( .B(n8979), .A(n8980), .S(n10649), .Y(n8978) );
  MUX2X1 U11436 ( .B(n8982), .A(n8983), .S(N21), .Y(n8981) );
  MUX2X1 U11437 ( .B(n8985), .A(n8986), .S(n10649), .Y(n8984) );
  MUX2X1 U11438 ( .B(n8988), .A(n8989), .S(n10649), .Y(n8987) );
  MUX2X1 U11439 ( .B(n8991), .A(n8992), .S(n10649), .Y(n8990) );
  MUX2X1 U11440 ( .B(n8994), .A(n8995), .S(n10649), .Y(n8993) );
  MUX2X1 U11441 ( .B(n8997), .A(n8998), .S(N21), .Y(n8996) );
  MUX2X1 U11442 ( .B(n9000), .A(n9001), .S(n10649), .Y(n8999) );
  MUX2X1 U11443 ( .B(n9003), .A(n9004), .S(n10649), .Y(n9002) );
  MUX2X1 U11444 ( .B(n9006), .A(n9007), .S(n10649), .Y(n9005) );
  MUX2X1 U11445 ( .B(n9009), .A(n9010), .S(n10649), .Y(n9008) );
  MUX2X1 U11446 ( .B(n9012), .A(n9013), .S(N21), .Y(n9011) );
  MUX2X1 U11447 ( .B(n9015), .A(n9016), .S(n10650), .Y(n9014) );
  MUX2X1 U11448 ( .B(n9018), .A(n9019), .S(n10650), .Y(n9017) );
  MUX2X1 U11449 ( .B(n9021), .A(n9022), .S(n10650), .Y(n9020) );
  MUX2X1 U11450 ( .B(n9024), .A(n9025), .S(n10650), .Y(n9023) );
  MUX2X1 U11451 ( .B(n9027), .A(n9028), .S(N21), .Y(n9026) );
  MUX2X1 U11452 ( .B(n9030), .A(n9031), .S(n10650), .Y(n9029) );
  MUX2X1 U11453 ( .B(n9033), .A(n9034), .S(n10650), .Y(n9032) );
  MUX2X1 U11454 ( .B(n9036), .A(n9037), .S(n10650), .Y(n9035) );
  MUX2X1 U11455 ( .B(n9039), .A(n9040), .S(n10650), .Y(n9038) );
  MUX2X1 U11456 ( .B(n9042), .A(n9043), .S(N21), .Y(n9041) );
  MUX2X1 U11457 ( .B(n9045), .A(n9046), .S(n10650), .Y(n9044) );
  MUX2X1 U11458 ( .B(n9048), .A(n9049), .S(n10650), .Y(n9047) );
  MUX2X1 U11459 ( .B(n9051), .A(n9052), .S(n10650), .Y(n9050) );
  MUX2X1 U11460 ( .B(n9054), .A(n9055), .S(n10650), .Y(n9053) );
  MUX2X1 U11461 ( .B(n9057), .A(n9058), .S(N21), .Y(n9056) );
  MUX2X1 U11462 ( .B(n9060), .A(n9061), .S(n10651), .Y(n9059) );
  MUX2X1 U11463 ( .B(n9063), .A(n9064), .S(n10651), .Y(n9062) );
  MUX2X1 U11464 ( .B(n9066), .A(n9067), .S(n10651), .Y(n9065) );
  MUX2X1 U11465 ( .B(n9069), .A(n9070), .S(n10651), .Y(n9068) );
  MUX2X1 U11466 ( .B(n9072), .A(n9073), .S(N21), .Y(n9071) );
  MUX2X1 U11467 ( .B(n9075), .A(n9076), .S(n10651), .Y(n9074) );
  MUX2X1 U11468 ( .B(n9078), .A(n9079), .S(n10651), .Y(n9077) );
  MUX2X1 U11469 ( .B(n9081), .A(n9082), .S(n10651), .Y(n9080) );
  MUX2X1 U11470 ( .B(n9084), .A(n9085), .S(n10651), .Y(n9083) );
  MUX2X1 U11471 ( .B(n9087), .A(n9088), .S(N21), .Y(n9086) );
  MUX2X1 U11472 ( .B(n9090), .A(n9091), .S(n10651), .Y(n9089) );
  MUX2X1 U11473 ( .B(n9093), .A(n9094), .S(n10651), .Y(n9092) );
  MUX2X1 U11474 ( .B(n9096), .A(n9097), .S(n10651), .Y(n9095) );
  MUX2X1 U11475 ( .B(n9099), .A(n9100), .S(n10651), .Y(n9098) );
  MUX2X1 U11476 ( .B(n9102), .A(n9103), .S(N21), .Y(n9101) );
  MUX2X1 U11477 ( .B(n9105), .A(n9106), .S(n10652), .Y(n9104) );
  MUX2X1 U11478 ( .B(n9108), .A(n9109), .S(n10652), .Y(n9107) );
  MUX2X1 U11479 ( .B(n9111), .A(n9112), .S(n10652), .Y(n9110) );
  MUX2X1 U11480 ( .B(n9114), .A(n9115), .S(n10652), .Y(n9113) );
  MUX2X1 U11481 ( .B(n9117), .A(n9118), .S(N21), .Y(n9116) );
  MUX2X1 U11482 ( .B(n9120), .A(n9121), .S(n10652), .Y(n9119) );
  MUX2X1 U11483 ( .B(n9123), .A(n9124), .S(n10652), .Y(n9122) );
  MUX2X1 U11484 ( .B(n9126), .A(n9127), .S(n10652), .Y(n9125) );
  MUX2X1 U11485 ( .B(n9129), .A(n9130), .S(n10652), .Y(n9128) );
  MUX2X1 U11486 ( .B(n9132), .A(n9133), .S(N21), .Y(n9131) );
  MUX2X1 U11487 ( .B(n9135), .A(n9136), .S(n10652), .Y(n9134) );
  MUX2X1 U11488 ( .B(n9138), .A(n9139), .S(n10652), .Y(n9137) );
  MUX2X1 U11489 ( .B(n9141), .A(n9142), .S(n10652), .Y(n9140) );
  MUX2X1 U11490 ( .B(n9144), .A(n9145), .S(n10652), .Y(n9143) );
  MUX2X1 U11491 ( .B(n9147), .A(n9148), .S(N21), .Y(n9146) );
  MUX2X1 U11492 ( .B(n9150), .A(n9151), .S(n10653), .Y(n9149) );
  MUX2X1 U11493 ( .B(n9153), .A(n9154), .S(n10653), .Y(n9152) );
  MUX2X1 U11494 ( .B(n9156), .A(n9157), .S(n10653), .Y(n9155) );
  MUX2X1 U11495 ( .B(n9159), .A(n9160), .S(n10653), .Y(n9158) );
  MUX2X1 U11496 ( .B(n9162), .A(n9163), .S(N21), .Y(n9161) );
  MUX2X1 U11497 ( .B(n9165), .A(n9166), .S(n10653), .Y(n9164) );
  MUX2X1 U11498 ( .B(n9168), .A(n9169), .S(n10653), .Y(n9167) );
  MUX2X1 U11499 ( .B(n9171), .A(n9172), .S(n10653), .Y(n9170) );
  MUX2X1 U11500 ( .B(n9174), .A(n9175), .S(n10653), .Y(n9173) );
  MUX2X1 U11501 ( .B(n9177), .A(n9178), .S(N21), .Y(n9176) );
  MUX2X1 U11502 ( .B(n9180), .A(n9181), .S(n10653), .Y(n9179) );
  MUX2X1 U11503 ( .B(n9183), .A(n9184), .S(n10653), .Y(n9182) );
  MUX2X1 U11504 ( .B(n9186), .A(n9187), .S(n10653), .Y(n9185) );
  MUX2X1 U11505 ( .B(n9189), .A(n9190), .S(n10653), .Y(n9188) );
  MUX2X1 U11506 ( .B(n9192), .A(n9193), .S(N21), .Y(n9191) );
  MUX2X1 U11507 ( .B(n9195), .A(n9196), .S(n10654), .Y(n9194) );
  MUX2X1 U11508 ( .B(n9198), .A(n9199), .S(n10654), .Y(n9197) );
  MUX2X1 U11509 ( .B(n9201), .A(n9202), .S(n10654), .Y(n9200) );
  MUX2X1 U11510 ( .B(n9204), .A(n9205), .S(n10654), .Y(n9203) );
  MUX2X1 U11511 ( .B(n9207), .A(n9208), .S(N21), .Y(n9206) );
  MUX2X1 U11512 ( .B(n9210), .A(n9211), .S(n10654), .Y(n9209) );
  MUX2X1 U11513 ( .B(n9213), .A(n9214), .S(n10654), .Y(n9212) );
  MUX2X1 U11514 ( .B(n9216), .A(n9217), .S(n10654), .Y(n9215) );
  MUX2X1 U11515 ( .B(n9219), .A(n9220), .S(n10654), .Y(n9218) );
  MUX2X1 U11516 ( .B(n9222), .A(n9223), .S(N21), .Y(n9221) );
  MUX2X1 U11517 ( .B(n9225), .A(n9226), .S(n10654), .Y(n9224) );
  MUX2X1 U11518 ( .B(n9228), .A(n9229), .S(n10654), .Y(n9227) );
  MUX2X1 U11519 ( .B(n9231), .A(n9232), .S(n10654), .Y(n9230) );
  MUX2X1 U11520 ( .B(n9234), .A(n9235), .S(n10654), .Y(n9233) );
  MUX2X1 U11521 ( .B(n9237), .A(n9238), .S(N21), .Y(n9236) );
  MUX2X1 U11522 ( .B(n9240), .A(n9241), .S(n10655), .Y(n9239) );
  MUX2X1 U11523 ( .B(n9243), .A(n9244), .S(n10655), .Y(n9242) );
  MUX2X1 U11524 ( .B(n9246), .A(n9247), .S(n10655), .Y(n9245) );
  MUX2X1 U11525 ( .B(n9249), .A(n9250), .S(n10655), .Y(n9248) );
  MUX2X1 U11526 ( .B(n9252), .A(n9253), .S(N21), .Y(n9251) );
  MUX2X1 U11527 ( .B(n9255), .A(n9256), .S(n10655), .Y(n9254) );
  MUX2X1 U11528 ( .B(n9258), .A(n9259), .S(n10655), .Y(n9257) );
  MUX2X1 U11529 ( .B(n9261), .A(n9262), .S(n10655), .Y(n9260) );
  MUX2X1 U11530 ( .B(n9264), .A(n9265), .S(n10655), .Y(n9263) );
  MUX2X1 U11531 ( .B(n9267), .A(n9268), .S(N21), .Y(n9266) );
  MUX2X1 U11532 ( .B(n9270), .A(n9271), .S(n10655), .Y(n9269) );
  MUX2X1 U11533 ( .B(n9273), .A(n9274), .S(n10655), .Y(n9272) );
  MUX2X1 U11534 ( .B(n9276), .A(n9277), .S(n10655), .Y(n9275) );
  MUX2X1 U11535 ( .B(n9279), .A(n9280), .S(n10655), .Y(n9278) );
  MUX2X1 U11536 ( .B(n9282), .A(n9283), .S(N21), .Y(n9281) );
  MUX2X1 U11537 ( .B(n9285), .A(n9286), .S(n10656), .Y(n9284) );
  MUX2X1 U11538 ( .B(n9288), .A(n9289), .S(n10656), .Y(n9287) );
  MUX2X1 U11539 ( .B(n9291), .A(n9292), .S(n10656), .Y(n9290) );
  MUX2X1 U11540 ( .B(n9294), .A(n9295), .S(n10656), .Y(n9293) );
  MUX2X1 U11541 ( .B(n9297), .A(n9298), .S(N21), .Y(n9296) );
  MUX2X1 U11542 ( .B(n9300), .A(n9301), .S(n10656), .Y(n9299) );
  MUX2X1 U11543 ( .B(n9303), .A(n9304), .S(n10656), .Y(n9302) );
  MUX2X1 U11544 ( .B(n9306), .A(n9307), .S(n10656), .Y(n9305) );
  MUX2X1 U11545 ( .B(n9309), .A(n9310), .S(n10656), .Y(n9308) );
  MUX2X1 U11546 ( .B(n9312), .A(n9313), .S(N21), .Y(n9311) );
  MUX2X1 U11547 ( .B(n9315), .A(n9316), .S(n10656), .Y(n9314) );
  MUX2X1 U11548 ( .B(n9318), .A(n9319), .S(n10656), .Y(n9317) );
  MUX2X1 U11549 ( .B(n9321), .A(n9322), .S(n10656), .Y(n9320) );
  MUX2X1 U11550 ( .B(n9324), .A(n9325), .S(n10656), .Y(n9323) );
  MUX2X1 U11551 ( .B(n9327), .A(n9328), .S(N21), .Y(n9326) );
  MUX2X1 U11552 ( .B(n9330), .A(n9331), .S(n10657), .Y(n9329) );
  MUX2X1 U11553 ( .B(n9333), .A(n9334), .S(n10657), .Y(n9332) );
  MUX2X1 U11554 ( .B(n9336), .A(n9337), .S(n10657), .Y(n9335) );
  MUX2X1 U11555 ( .B(n9339), .A(n9340), .S(n10657), .Y(n9338) );
  MUX2X1 U11556 ( .B(n9342), .A(n9343), .S(N21), .Y(n9341) );
  MUX2X1 U11557 ( .B(n9345), .A(n9346), .S(n10657), .Y(n9344) );
  MUX2X1 U11558 ( .B(n9348), .A(n9349), .S(n10657), .Y(n9347) );
  MUX2X1 U11559 ( .B(n9351), .A(n9352), .S(n10657), .Y(n9350) );
  MUX2X1 U11560 ( .B(n9354), .A(n9355), .S(n10657), .Y(n9353) );
  MUX2X1 U11561 ( .B(n9357), .A(n9358), .S(N21), .Y(n9356) );
  MUX2X1 U11562 ( .B(n9360), .A(n9361), .S(n10657), .Y(n9359) );
  MUX2X1 U11563 ( .B(n9363), .A(n9364), .S(n10657), .Y(n9362) );
  MUX2X1 U11564 ( .B(n9366), .A(n9367), .S(n10657), .Y(n9365) );
  MUX2X1 U11565 ( .B(n9369), .A(n9370), .S(n10657), .Y(n9368) );
  MUX2X1 U11566 ( .B(n9372), .A(n9373), .S(N21), .Y(n9371) );
  MUX2X1 U11567 ( .B(n9375), .A(n9376), .S(n10658), .Y(n9374) );
  MUX2X1 U11568 ( .B(n9378), .A(n9379), .S(n10658), .Y(n9377) );
  MUX2X1 U11569 ( .B(n9381), .A(n9382), .S(n10658), .Y(n9380) );
  MUX2X1 U11570 ( .B(n9384), .A(n9385), .S(n10658), .Y(n9383) );
  MUX2X1 U11571 ( .B(n9387), .A(n9388), .S(N21), .Y(n9386) );
  MUX2X1 U11572 ( .B(n9390), .A(n9391), .S(n10658), .Y(n9389) );
  MUX2X1 U11573 ( .B(n9393), .A(n9394), .S(n10658), .Y(n9392) );
  MUX2X1 U11574 ( .B(n9396), .A(n9397), .S(n10658), .Y(n9395) );
  MUX2X1 U11575 ( .B(n9399), .A(n9400), .S(n10658), .Y(n9398) );
  MUX2X1 U11576 ( .B(n9402), .A(n9403), .S(N21), .Y(n9401) );
  MUX2X1 U11577 ( .B(n9405), .A(n9406), .S(n10658), .Y(n9404) );
  MUX2X1 U11578 ( .B(n9408), .A(n9409), .S(n10658), .Y(n9407) );
  MUX2X1 U11579 ( .B(n9411), .A(n9412), .S(n10658), .Y(n9410) );
  MUX2X1 U11580 ( .B(n9414), .A(n9415), .S(n10658), .Y(n9413) );
  MUX2X1 U11581 ( .B(n9417), .A(n9418), .S(N21), .Y(n9416) );
  MUX2X1 U11582 ( .B(n9420), .A(n9421), .S(n10659), .Y(n9419) );
  MUX2X1 U11583 ( .B(n9423), .A(n9424), .S(n10659), .Y(n9422) );
  MUX2X1 U11584 ( .B(n9426), .A(n9427), .S(n10659), .Y(n9425) );
  MUX2X1 U11585 ( .B(n9429), .A(n9430), .S(n10659), .Y(n9428) );
  MUX2X1 U11586 ( .B(n9432), .A(n9433), .S(N21), .Y(n9431) );
  MUX2X1 U11587 ( .B(n9435), .A(n9436), .S(n10659), .Y(n9434) );
  MUX2X1 U11588 ( .B(n9438), .A(n9439), .S(n10659), .Y(n9437) );
  MUX2X1 U11589 ( .B(n9441), .A(n9442), .S(n10659), .Y(n9440) );
  MUX2X1 U11590 ( .B(n9444), .A(n9445), .S(n10659), .Y(n9443) );
  MUX2X1 U11591 ( .B(n9447), .A(n9448), .S(N21), .Y(n9446) );
  MUX2X1 U11592 ( .B(n9450), .A(n9451), .S(n10659), .Y(n9449) );
  MUX2X1 U11593 ( .B(n9453), .A(n9454), .S(n10659), .Y(n9452) );
  MUX2X1 U11594 ( .B(n9456), .A(n9457), .S(n10659), .Y(n9455) );
  MUX2X1 U11595 ( .B(n9459), .A(n9460), .S(n10659), .Y(n9458) );
  MUX2X1 U11596 ( .B(n9462), .A(n9463), .S(N21), .Y(n9461) );
  MUX2X1 U11597 ( .B(n9465), .A(n9466), .S(n10660), .Y(n9464) );
  MUX2X1 U11598 ( .B(n9468), .A(n9469), .S(n10660), .Y(n9467) );
  MUX2X1 U11599 ( .B(n9471), .A(n9472), .S(n10660), .Y(n9470) );
  MUX2X1 U11600 ( .B(n9474), .A(n9475), .S(n10660), .Y(n9473) );
  MUX2X1 U11601 ( .B(n9477), .A(n9478), .S(N21), .Y(n9476) );
  MUX2X1 U11602 ( .B(n9480), .A(n9481), .S(n10660), .Y(n9479) );
  MUX2X1 U11603 ( .B(n9483), .A(n9484), .S(n10660), .Y(n9482) );
  MUX2X1 U11604 ( .B(n9486), .A(n9487), .S(n10660), .Y(n9485) );
  MUX2X1 U11605 ( .B(n9489), .A(n9490), .S(n10660), .Y(n9488) );
  MUX2X1 U11606 ( .B(n9492), .A(n9493), .S(N21), .Y(n9491) );
  MUX2X1 U11607 ( .B(n9495), .A(n9496), .S(n10660), .Y(n9494) );
  MUX2X1 U11608 ( .B(n9498), .A(n9499), .S(n10660), .Y(n9497) );
  MUX2X1 U11609 ( .B(n9501), .A(n9502), .S(n10660), .Y(n9500) );
  MUX2X1 U11610 ( .B(n9504), .A(n9505), .S(n10660), .Y(n9503) );
  MUX2X1 U11611 ( .B(n9507), .A(n9508), .S(N21), .Y(n9506) );
  MUX2X1 U11612 ( .B(n9510), .A(n9511), .S(n10661), .Y(n9509) );
  MUX2X1 U11613 ( .B(n9513), .A(n9514), .S(n10661), .Y(n9512) );
  MUX2X1 U11614 ( .B(n9516), .A(n9517), .S(n10661), .Y(n9515) );
  MUX2X1 U11615 ( .B(n9519), .A(n9520), .S(n10661), .Y(n9518) );
  MUX2X1 U11616 ( .B(n9522), .A(n9523), .S(N21), .Y(n9521) );
  MUX2X1 U11617 ( .B(n9525), .A(n9526), .S(n10661), .Y(n9524) );
  MUX2X1 U11618 ( .B(n9528), .A(n9529), .S(n10661), .Y(n9527) );
  MUX2X1 U11619 ( .B(n9531), .A(n9532), .S(n10661), .Y(n9530) );
  MUX2X1 U11620 ( .B(n9534), .A(n9535), .S(n10661), .Y(n9533) );
  MUX2X1 U11621 ( .B(n9537), .A(n9538), .S(N21), .Y(n9536) );
  MUX2X1 U11622 ( .B(n9540), .A(n9541), .S(n10661), .Y(n9539) );
  MUX2X1 U11623 ( .B(n9543), .A(n9544), .S(n10661), .Y(n9542) );
  MUX2X1 U11624 ( .B(n9546), .A(n9547), .S(n10661), .Y(n9545) );
  MUX2X1 U11625 ( .B(n9549), .A(n9550), .S(n10661), .Y(n9548) );
  MUX2X1 U11626 ( .B(n9552), .A(n9553), .S(N21), .Y(n9551) );
  MUX2X1 U11627 ( .B(n9555), .A(n9556), .S(n10662), .Y(n9554) );
  MUX2X1 U11628 ( .B(n9558), .A(n9559), .S(n10662), .Y(n9557) );
  MUX2X1 U11629 ( .B(n9561), .A(n9562), .S(n10662), .Y(n9560) );
  MUX2X1 U11630 ( .B(n9564), .A(n9565), .S(n10662), .Y(n9563) );
  MUX2X1 U11631 ( .B(n9567), .A(n9568), .S(N21), .Y(n9566) );
  MUX2X1 U11632 ( .B(n9570), .A(n9571), .S(n10662), .Y(n9569) );
  MUX2X1 U11633 ( .B(n9573), .A(n9574), .S(n10662), .Y(n9572) );
  MUX2X1 U11634 ( .B(n9576), .A(n9577), .S(n10662), .Y(n9575) );
  MUX2X1 U11635 ( .B(n9579), .A(n9580), .S(n10662), .Y(n9578) );
  MUX2X1 U11636 ( .B(n9582), .A(n9583), .S(N21), .Y(n9581) );
  MUX2X1 U11637 ( .B(n9585), .A(n9586), .S(n10662), .Y(n9584) );
  MUX2X1 U11638 ( .B(n9588), .A(n9589), .S(n10662), .Y(n9587) );
  MUX2X1 U11639 ( .B(n9591), .A(n9592), .S(n10662), .Y(n9590) );
  MUX2X1 U11640 ( .B(n9594), .A(n9595), .S(n10662), .Y(n9593) );
  MUX2X1 U11641 ( .B(n9597), .A(n9598), .S(N21), .Y(n9596) );
  MUX2X1 U11642 ( .B(n9600), .A(n9601), .S(n10663), .Y(n9599) );
  MUX2X1 U11643 ( .B(n9603), .A(n9604), .S(n10663), .Y(n9602) );
  MUX2X1 U11644 ( .B(n9606), .A(n9607), .S(n10663), .Y(n9605) );
  MUX2X1 U11645 ( .B(n9609), .A(n9610), .S(n10663), .Y(n9608) );
  MUX2X1 U11646 ( .B(n9612), .A(n9613), .S(N21), .Y(n9611) );
  MUX2X1 U11647 ( .B(n9615), .A(n9616), .S(n10663), .Y(n9614) );
  MUX2X1 U11648 ( .B(n9618), .A(n9619), .S(n10663), .Y(n9617) );
  MUX2X1 U11649 ( .B(n9621), .A(n9622), .S(n10663), .Y(n9620) );
  MUX2X1 U11650 ( .B(n9624), .A(n9625), .S(n10663), .Y(n9623) );
  MUX2X1 U11651 ( .B(n9627), .A(n9628), .S(N21), .Y(n9626) );
  MUX2X1 U11652 ( .B(n9630), .A(n9631), .S(n10663), .Y(n9629) );
  MUX2X1 U11653 ( .B(n9633), .A(n9634), .S(n10663), .Y(n9632) );
  MUX2X1 U11654 ( .B(n9636), .A(n9637), .S(n10663), .Y(n9635) );
  MUX2X1 U11655 ( .B(n9639), .A(n9640), .S(n10663), .Y(n9638) );
  MUX2X1 U11656 ( .B(n9642), .A(n9643), .S(N21), .Y(n9641) );
  MUX2X1 U11657 ( .B(n9645), .A(n9646), .S(n10664), .Y(n9644) );
  MUX2X1 U11658 ( .B(n9648), .A(n9649), .S(n10664), .Y(n9647) );
  MUX2X1 U11659 ( .B(n9651), .A(n9652), .S(n10664), .Y(n9650) );
  MUX2X1 U11660 ( .B(n9654), .A(n9655), .S(n10664), .Y(n9653) );
  MUX2X1 U11661 ( .B(n9657), .A(n9658), .S(N21), .Y(n9656) );
  MUX2X1 U11662 ( .B(n9660), .A(n9661), .S(n10664), .Y(n9659) );
  MUX2X1 U11663 ( .B(n9663), .A(n9664), .S(n10664), .Y(n9662) );
  MUX2X1 U11664 ( .B(n9666), .A(n9667), .S(n10664), .Y(n9665) );
  MUX2X1 U11665 ( .B(n9669), .A(n9670), .S(n10664), .Y(n9668) );
  MUX2X1 U11666 ( .B(n9672), .A(n9673), .S(N21), .Y(n9671) );
  MUX2X1 U11667 ( .B(n9675), .A(n9676), .S(n10664), .Y(n9674) );
  MUX2X1 U11668 ( .B(n9678), .A(n9679), .S(n10664), .Y(n9677) );
  MUX2X1 U11669 ( .B(n9681), .A(n9682), .S(n10664), .Y(n9680) );
  MUX2X1 U11670 ( .B(n9684), .A(n9685), .S(n10664), .Y(n9683) );
  MUX2X1 U11671 ( .B(n9687), .A(n9688), .S(N21), .Y(n9686) );
  MUX2X1 U11672 ( .B(n9690), .A(n9691), .S(n10665), .Y(n9689) );
  MUX2X1 U11673 ( .B(n9693), .A(n9694), .S(n10665), .Y(n9692) );
  MUX2X1 U11674 ( .B(n9696), .A(n9697), .S(n10665), .Y(n9695) );
  MUX2X1 U11675 ( .B(n9699), .A(n9700), .S(n10665), .Y(n9698) );
  MUX2X1 U11676 ( .B(n9702), .A(n9703), .S(N21), .Y(n9701) );
  MUX2X1 U11677 ( .B(n9705), .A(n9706), .S(n10665), .Y(n9704) );
  MUX2X1 U11678 ( .B(n9708), .A(n9709), .S(n10665), .Y(n9707) );
  MUX2X1 U11679 ( .B(n9711), .A(n9712), .S(n10665), .Y(n9710) );
  MUX2X1 U11680 ( .B(n9714), .A(n9715), .S(n10665), .Y(n9713) );
  MUX2X1 U11681 ( .B(n9717), .A(n9718), .S(N21), .Y(n9716) );
  MUX2X1 U11682 ( .B(n9720), .A(n9721), .S(n10665), .Y(n9719) );
  MUX2X1 U11683 ( .B(n9723), .A(n9724), .S(n10665), .Y(n9722) );
  MUX2X1 U11684 ( .B(n9726), .A(n9727), .S(n10665), .Y(n9725) );
  MUX2X1 U11685 ( .B(n9729), .A(n9730), .S(n10665), .Y(n9728) );
  MUX2X1 U11686 ( .B(n9732), .A(n9733), .S(N21), .Y(n9731) );
  MUX2X1 U11687 ( .B(n9735), .A(n9736), .S(n10666), .Y(n9734) );
  MUX2X1 U11688 ( .B(n9738), .A(n9739), .S(n10666), .Y(n9737) );
  MUX2X1 U11689 ( .B(n9741), .A(n9742), .S(n10666), .Y(n9740) );
  MUX2X1 U11690 ( .B(n9744), .A(n9745), .S(n10666), .Y(n9743) );
  MUX2X1 U11691 ( .B(n9747), .A(n9748), .S(N21), .Y(n9746) );
  MUX2X1 U11692 ( .B(n9750), .A(n9751), .S(n10666), .Y(n9749) );
  MUX2X1 U11693 ( .B(n9753), .A(n9754), .S(n10666), .Y(n9752) );
  MUX2X1 U11694 ( .B(n9756), .A(n9757), .S(n10666), .Y(n9755) );
  MUX2X1 U11695 ( .B(n9759), .A(n9760), .S(n10666), .Y(n9758) );
  MUX2X1 U11696 ( .B(n9762), .A(n9763), .S(N21), .Y(n9761) );
  MUX2X1 U11697 ( .B(n9765), .A(n9766), .S(n10666), .Y(n9764) );
  MUX2X1 U11698 ( .B(n9768), .A(n9769), .S(n10666), .Y(n9767) );
  MUX2X1 U11699 ( .B(n9771), .A(n9772), .S(n10666), .Y(n9770) );
  MUX2X1 U11700 ( .B(n9774), .A(n9775), .S(n10666), .Y(n9773) );
  MUX2X1 U11701 ( .B(n9777), .A(n9778), .S(N21), .Y(n9776) );
  MUX2X1 U11702 ( .B(n9780), .A(n9781), .S(n10667), .Y(n9779) );
  MUX2X1 U11703 ( .B(n9783), .A(n9784), .S(n10667), .Y(n9782) );
  MUX2X1 U11704 ( .B(n9786), .A(n9787), .S(n10667), .Y(n9785) );
  MUX2X1 U11705 ( .B(n9789), .A(n9790), .S(n10667), .Y(n9788) );
  MUX2X1 U11706 ( .B(n9792), .A(n9793), .S(N21), .Y(n9791) );
  MUX2X1 U11707 ( .B(n9795), .A(n9796), .S(n10667), .Y(n9794) );
  MUX2X1 U11708 ( .B(n9798), .A(n9799), .S(n10667), .Y(n9797) );
  MUX2X1 U11709 ( .B(n9801), .A(n9802), .S(n10667), .Y(n9800) );
  MUX2X1 U11710 ( .B(n9804), .A(n9805), .S(n10667), .Y(n9803) );
  MUX2X1 U11711 ( .B(n9807), .A(n9808), .S(N21), .Y(n9806) );
  MUX2X1 U11712 ( .B(n9810), .A(n9811), .S(n10667), .Y(n9809) );
  MUX2X1 U11713 ( .B(n9813), .A(n9814), .S(n10667), .Y(n9812) );
  MUX2X1 U11714 ( .B(n9816), .A(n9817), .S(n10667), .Y(n9815) );
  MUX2X1 U11715 ( .B(n9819), .A(n9820), .S(n10667), .Y(n9818) );
  MUX2X1 U11716 ( .B(n9822), .A(n9823), .S(N21), .Y(n9821) );
  MUX2X1 U11717 ( .B(n9825), .A(n9826), .S(n10668), .Y(n9824) );
  MUX2X1 U11718 ( .B(n9828), .A(n9829), .S(n10668), .Y(n9827) );
  MUX2X1 U11719 ( .B(n9831), .A(n9832), .S(n10668), .Y(n9830) );
  MUX2X1 U11720 ( .B(n9834), .A(n9835), .S(n10668), .Y(n9833) );
  MUX2X1 U11721 ( .B(n9837), .A(n9838), .S(N21), .Y(n9836) );
  MUX2X1 U11722 ( .B(n9840), .A(n9841), .S(n10668), .Y(n9839) );
  MUX2X1 U11723 ( .B(n9843), .A(n9844), .S(n10668), .Y(n9842) );
  MUX2X1 U11724 ( .B(n9846), .A(n9847), .S(n10668), .Y(n9845) );
  MUX2X1 U11725 ( .B(n9849), .A(n9850), .S(n10668), .Y(n9848) );
  MUX2X1 U11726 ( .B(n9852), .A(n9853), .S(N21), .Y(n9851) );
  MUX2X1 U11727 ( .B(n9855), .A(n9856), .S(n10668), .Y(n9854) );
  MUX2X1 U11728 ( .B(n9858), .A(n9859), .S(n10668), .Y(n9857) );
  MUX2X1 U11729 ( .B(n9861), .A(n9862), .S(n10668), .Y(n9860) );
  MUX2X1 U11730 ( .B(n9864), .A(n9865), .S(n10668), .Y(n9863) );
  MUX2X1 U11731 ( .B(n9867), .A(n9868), .S(N21), .Y(n9866) );
  MUX2X1 U11732 ( .B(n9870), .A(n9871), .S(n10669), .Y(n9869) );
  MUX2X1 U11733 ( .B(n9873), .A(n9874), .S(n10669), .Y(n9872) );
  MUX2X1 U11734 ( .B(n9876), .A(n9877), .S(n10669), .Y(n9875) );
  MUX2X1 U11735 ( .B(n9879), .A(n9880), .S(n10669), .Y(n9878) );
  MUX2X1 U11736 ( .B(n9882), .A(n9883), .S(N21), .Y(n9881) );
  MUX2X1 U11737 ( .B(n9885), .A(n9886), .S(n10669), .Y(n9884) );
  MUX2X1 U11738 ( .B(n9888), .A(n9889), .S(n10669), .Y(n9887) );
  MUX2X1 U11739 ( .B(n9891), .A(n9892), .S(n10669), .Y(n9890) );
  MUX2X1 U11740 ( .B(n9894), .A(n9895), .S(n10669), .Y(n9893) );
  MUX2X1 U11741 ( .B(n9897), .A(n9898), .S(N21), .Y(n9896) );
  MUX2X1 U11742 ( .B(n9900), .A(n9901), .S(n10669), .Y(n9899) );
  MUX2X1 U11743 ( .B(n9903), .A(n9904), .S(n10669), .Y(n9902) );
  MUX2X1 U11744 ( .B(n9906), .A(n9907), .S(n10669), .Y(n9905) );
  MUX2X1 U11745 ( .B(n9909), .A(n9910), .S(n10669), .Y(n9908) );
  MUX2X1 U11746 ( .B(n9912), .A(n9913), .S(N21), .Y(n9911) );
  MUX2X1 U11747 ( .B(n9915), .A(n9916), .S(n10670), .Y(n9914) );
  MUX2X1 U11748 ( .B(n9918), .A(n9919), .S(n10670), .Y(n9917) );
  MUX2X1 U11749 ( .B(n9921), .A(n9922), .S(n10670), .Y(n9920) );
  MUX2X1 U11750 ( .B(n9924), .A(n9925), .S(n10670), .Y(n9923) );
  MUX2X1 U11751 ( .B(n9927), .A(n9928), .S(N21), .Y(n9926) );
  MUX2X1 U11752 ( .B(n9930), .A(n9931), .S(n10670), .Y(n9929) );
  MUX2X1 U11753 ( .B(n9933), .A(n9934), .S(n10670), .Y(n9932) );
  MUX2X1 U11754 ( .B(n9936), .A(n9937), .S(n10670), .Y(n9935) );
  MUX2X1 U11755 ( .B(n9939), .A(n9940), .S(n10670), .Y(n9938) );
  MUX2X1 U11756 ( .B(n9942), .A(n9943), .S(N21), .Y(n9941) );
  MUX2X1 U11757 ( .B(n9945), .A(n9946), .S(n10670), .Y(n9944) );
  MUX2X1 U11758 ( .B(n9948), .A(n9949), .S(n10670), .Y(n9947) );
  MUX2X1 U11759 ( .B(n9951), .A(n9952), .S(n10670), .Y(n9950) );
  MUX2X1 U11760 ( .B(n9954), .A(n9955), .S(n10670), .Y(n9953) );
  MUX2X1 U11761 ( .B(n9957), .A(n9958), .S(N21), .Y(n9956) );
  MUX2X1 U11762 ( .B(n9960), .A(n9961), .S(n10671), .Y(n9959) );
  MUX2X1 U11763 ( .B(n9963), .A(n9964), .S(n10671), .Y(n9962) );
  MUX2X1 U11764 ( .B(n9966), .A(n9967), .S(n10671), .Y(n9965) );
  MUX2X1 U11765 ( .B(n9969), .A(n9970), .S(n10671), .Y(n9968) );
  MUX2X1 U11766 ( .B(n9972), .A(n9973), .S(N21), .Y(n9971) );
  MUX2X1 U11767 ( .B(n9975), .A(n9976), .S(n10671), .Y(n9974) );
  MUX2X1 U11768 ( .B(n9978), .A(n9979), .S(n10671), .Y(n9977) );
  MUX2X1 U11769 ( .B(n9981), .A(n9982), .S(n10671), .Y(n9980) );
  MUX2X1 U11770 ( .B(n9984), .A(n9985), .S(n10671), .Y(n9983) );
  MUX2X1 U11771 ( .B(n9987), .A(n9988), .S(N21), .Y(n9986) );
  MUX2X1 U11772 ( .B(n9990), .A(n9991), .S(n10671), .Y(n9989) );
  MUX2X1 U11773 ( .B(n9993), .A(n9994), .S(n10671), .Y(n9992) );
  MUX2X1 U11774 ( .B(n9996), .A(n9997), .S(n10671), .Y(n9995) );
  MUX2X1 U11775 ( .B(n9999), .A(n10000), .S(n10671), .Y(n9998) );
  MUX2X1 U11776 ( .B(n10002), .A(n10003), .S(N21), .Y(n10001) );
  MUX2X1 U11777 ( .B(n10005), .A(n10006), .S(n10672), .Y(n10004) );
  MUX2X1 U11778 ( .B(n10008), .A(n10009), .S(n10672), .Y(n10007) );
  MUX2X1 U11779 ( .B(n10011), .A(n10012), .S(n10672), .Y(n10010) );
  MUX2X1 U11780 ( .B(n10014), .A(n10015), .S(n10672), .Y(n10013) );
  MUX2X1 U11781 ( .B(n10017), .A(n10018), .S(N21), .Y(n10016) );
  MUX2X1 U11782 ( .B(n10020), .A(n10021), .S(n10672), .Y(n10019) );
  MUX2X1 U11783 ( .B(n10023), .A(n10024), .S(n10672), .Y(n10022) );
  MUX2X1 U11784 ( .B(n10026), .A(n10027), .S(n10672), .Y(n10025) );
  MUX2X1 U11785 ( .B(n10029), .A(n10030), .S(n10672), .Y(n10028) );
  MUX2X1 U11786 ( .B(n10032), .A(n10033), .S(N21), .Y(n10031) );
  MUX2X1 U11787 ( .B(n10035), .A(n10036), .S(n10672), .Y(n10034) );
  MUX2X1 U11788 ( .B(n10038), .A(n10039), .S(n10672), .Y(n10037) );
  MUX2X1 U11789 ( .B(n10041), .A(n10042), .S(n10672), .Y(n10040) );
  MUX2X1 U11790 ( .B(n10044), .A(n10045), .S(n10672), .Y(n10043) );
  MUX2X1 U11791 ( .B(n10047), .A(n10048), .S(N21), .Y(n10046) );
  MUX2X1 U11792 ( .B(n10050), .A(n10051), .S(n10673), .Y(n10049) );
  MUX2X1 U11793 ( .B(n10053), .A(n10054), .S(n10673), .Y(n10052) );
  MUX2X1 U11794 ( .B(n10056), .A(n10057), .S(n10673), .Y(n10055) );
  MUX2X1 U11795 ( .B(n10059), .A(n10060), .S(n10673), .Y(n10058) );
  MUX2X1 U11796 ( .B(n10062), .A(n10063), .S(N21), .Y(n10061) );
  MUX2X1 U11797 ( .B(n10065), .A(n10066), .S(n10673), .Y(n10064) );
  MUX2X1 U11798 ( .B(n10068), .A(n10069), .S(n10673), .Y(n10067) );
  MUX2X1 U11799 ( .B(n10071), .A(n10072), .S(n10673), .Y(n10070) );
  MUX2X1 U11800 ( .B(n10074), .A(n10075), .S(n10673), .Y(n10073) );
  MUX2X1 U11801 ( .B(n10077), .A(n10078), .S(N21), .Y(n10076) );
  MUX2X1 U11802 ( .B(n10080), .A(n10081), .S(n10673), .Y(n10079) );
  MUX2X1 U11803 ( .B(n10083), .A(n10084), .S(n10673), .Y(n10082) );
  MUX2X1 U11804 ( .B(n10086), .A(n10087), .S(n10673), .Y(n10085) );
  MUX2X1 U11805 ( .B(n10089), .A(n10090), .S(n10673), .Y(n10088) );
  MUX2X1 U11806 ( .B(n10092), .A(n10093), .S(N21), .Y(n10091) );
  MUX2X1 U11807 ( .B(n10095), .A(n10096), .S(n10674), .Y(n10094) );
  MUX2X1 U11808 ( .B(n10098), .A(n10099), .S(n10674), .Y(n10097) );
  MUX2X1 U11809 ( .B(n10101), .A(n10102), .S(n10674), .Y(n10100) );
  MUX2X1 U11810 ( .B(n10104), .A(n10105), .S(n10674), .Y(n10103) );
  MUX2X1 U11811 ( .B(n10107), .A(n10108), .S(N21), .Y(n10106) );
  MUX2X1 U11812 ( .B(n10110), .A(n10111), .S(n10674), .Y(n10109) );
  MUX2X1 U11813 ( .B(n10113), .A(n10114), .S(n10674), .Y(n10112) );
  MUX2X1 U11814 ( .B(n10116), .A(n10117), .S(n10674), .Y(n10115) );
  MUX2X1 U11815 ( .B(n10119), .A(n10120), .S(n10674), .Y(n10118) );
  MUX2X1 U11816 ( .B(n10122), .A(n10123), .S(N21), .Y(n10121) );
  MUX2X1 U11817 ( .B(n10125), .A(n10126), .S(n10674), .Y(n10124) );
  MUX2X1 U11818 ( .B(n10128), .A(n10129), .S(n10674), .Y(n10127) );
  MUX2X1 U11819 ( .B(n10131), .A(n10132), .S(n10674), .Y(n10130) );
  MUX2X1 U11820 ( .B(n10134), .A(n10135), .S(n10674), .Y(n10133) );
  MUX2X1 U11821 ( .B(n10137), .A(n10138), .S(N21), .Y(n10136) );
  MUX2X1 U11822 ( .B(n10140), .A(n10141), .S(n10675), .Y(n10139) );
  MUX2X1 U11823 ( .B(n10143), .A(n10144), .S(n10675), .Y(n10142) );
  MUX2X1 U11824 ( .B(n10146), .A(n10147), .S(n10675), .Y(n10145) );
  MUX2X1 U11825 ( .B(n10149), .A(n10150), .S(n10675), .Y(n10148) );
  MUX2X1 U11826 ( .B(n10152), .A(n10153), .S(N21), .Y(n10151) );
  MUX2X1 U11827 ( .B(n10155), .A(n10156), .S(n10675), .Y(n10154) );
  MUX2X1 U11828 ( .B(n10158), .A(n10159), .S(n10675), .Y(n10157) );
  MUX2X1 U11829 ( .B(n10161), .A(n10162), .S(n10675), .Y(n10160) );
  MUX2X1 U11830 ( .B(n10164), .A(n10165), .S(n10675), .Y(n10163) );
  MUX2X1 U11831 ( .B(n10167), .A(n10168), .S(N21), .Y(n10166) );
  MUX2X1 U11832 ( .B(n10170), .A(n10171), .S(n10675), .Y(n10169) );
  MUX2X1 U11833 ( .B(n10173), .A(n10174), .S(n10675), .Y(n10172) );
  MUX2X1 U11834 ( .B(n10176), .A(n10177), .S(n10675), .Y(n10175) );
  MUX2X1 U11835 ( .B(n10179), .A(n10180), .S(n10675), .Y(n10178) );
  MUX2X1 U11836 ( .B(n10182), .A(n10183), .S(N21), .Y(n10181) );
  MUX2X1 U11837 ( .B(n10185), .A(n10186), .S(n10676), .Y(n10184) );
  MUX2X1 U11838 ( .B(n10188), .A(n10189), .S(n10676), .Y(n10187) );
  MUX2X1 U11839 ( .B(n10191), .A(n10192), .S(n10676), .Y(n10190) );
  MUX2X1 U11840 ( .B(n10194), .A(n10195), .S(n10676), .Y(n10193) );
  MUX2X1 U11841 ( .B(n10197), .A(n10198), .S(N21), .Y(n10196) );
  MUX2X1 U11842 ( .B(n10200), .A(n10201), .S(n10676), .Y(n10199) );
  MUX2X1 U11843 ( .B(n10203), .A(n10204), .S(n10676), .Y(n10202) );
  MUX2X1 U11844 ( .B(n10206), .A(n10207), .S(n10676), .Y(n10205) );
  MUX2X1 U11845 ( .B(n10209), .A(n10210), .S(n10676), .Y(n10208) );
  MUX2X1 U11846 ( .B(n10212), .A(n10213), .S(N21), .Y(n10211) );
  MUX2X1 U11847 ( .B(n10215), .A(n10216), .S(n10676), .Y(n10214) );
  MUX2X1 U11848 ( .B(n10218), .A(n10219), .S(n10676), .Y(n10217) );
  MUX2X1 U11849 ( .B(n10221), .A(n10222), .S(n10676), .Y(n10220) );
  MUX2X1 U11850 ( .B(n10224), .A(n10225), .S(n10676), .Y(n10223) );
  MUX2X1 U11851 ( .B(n10227), .A(n10228), .S(N21), .Y(n10226) );
  MUX2X1 U11852 ( .B(n10230), .A(n10231), .S(n10677), .Y(n10229) );
  MUX2X1 U11853 ( .B(n10233), .A(n10234), .S(n10677), .Y(n10232) );
  MUX2X1 U11854 ( .B(n10236), .A(n10237), .S(n10677), .Y(n10235) );
  MUX2X1 U11855 ( .B(n10239), .A(n10240), .S(n10677), .Y(n10238) );
  MUX2X1 U11856 ( .B(n10242), .A(n10243), .S(N21), .Y(n10241) );
  MUX2X1 U11857 ( .B(n10245), .A(n10246), .S(n10677), .Y(n10244) );
  MUX2X1 U11858 ( .B(n10248), .A(n10249), .S(n10677), .Y(n10247) );
  MUX2X1 U11859 ( .B(n10251), .A(n10252), .S(n10677), .Y(n10250) );
  MUX2X1 U11860 ( .B(n10254), .A(n10255), .S(n10677), .Y(n10253) );
  MUX2X1 U11861 ( .B(n10257), .A(n10258), .S(N21), .Y(n10256) );
  MUX2X1 U11862 ( .B(n10260), .A(n10261), .S(n10677), .Y(n10259) );
  MUX2X1 U11863 ( .B(n10263), .A(n10264), .S(n10677), .Y(n10262) );
  MUX2X1 U11864 ( .B(n10266), .A(n10267), .S(n10677), .Y(n10265) );
  MUX2X1 U11865 ( .B(n10269), .A(n10270), .S(n10677), .Y(n10268) );
  MUX2X1 U11866 ( .B(n10272), .A(n10273), .S(N21), .Y(n10271) );
  MUX2X1 U11867 ( .B(n10275), .A(n10276), .S(n10678), .Y(n10274) );
  MUX2X1 U11868 ( .B(n10278), .A(n10279), .S(n10678), .Y(n10277) );
  MUX2X1 U11869 ( .B(n10281), .A(n10282), .S(n10678), .Y(n10280) );
  MUX2X1 U11870 ( .B(n10284), .A(n10285), .S(n10678), .Y(n10283) );
  MUX2X1 U11871 ( .B(n10287), .A(n10288), .S(N21), .Y(n10286) );
  MUX2X1 U11872 ( .B(n10290), .A(n10291), .S(n10678), .Y(n10289) );
  MUX2X1 U11873 ( .B(n10293), .A(n10294), .S(n10678), .Y(n10292) );
  MUX2X1 U11874 ( .B(n10296), .A(n10297), .S(n10678), .Y(n10295) );
  MUX2X1 U11875 ( .B(n10299), .A(n10300), .S(n10678), .Y(n10298) );
  MUX2X1 U11876 ( .B(n10302), .A(n10303), .S(N21), .Y(n10301) );
  MUX2X1 U11877 ( .B(n10305), .A(n10306), .S(n10678), .Y(n10304) );
  MUX2X1 U11878 ( .B(n10308), .A(n10309), .S(n10678), .Y(n10307) );
  MUX2X1 U11879 ( .B(n10311), .A(n10312), .S(n10678), .Y(n10310) );
  MUX2X1 U11880 ( .B(n10314), .A(n10315), .S(n10678), .Y(n10313) );
  MUX2X1 U11881 ( .B(n10317), .A(n10318), .S(N21), .Y(n10316) );
  MUX2X1 U11882 ( .B(n10320), .A(n10321), .S(n10679), .Y(n10319) );
  MUX2X1 U11883 ( .B(n10323), .A(n10324), .S(n10679), .Y(n10322) );
  MUX2X1 U11884 ( .B(n10326), .A(n10327), .S(n10679), .Y(n10325) );
  MUX2X1 U11885 ( .B(n10329), .A(n10330), .S(n10679), .Y(n10328) );
  MUX2X1 U11886 ( .B(n10332), .A(n10333), .S(N21), .Y(n10331) );
  MUX2X1 U11887 ( .B(n10335), .A(n10336), .S(n10679), .Y(n10334) );
  MUX2X1 U11888 ( .B(n10338), .A(n10339), .S(n10679), .Y(n10337) );
  MUX2X1 U11889 ( .B(n10341), .A(n10342), .S(n10679), .Y(n10340) );
  MUX2X1 U11890 ( .B(n10344), .A(n10345), .S(n10679), .Y(n10343) );
  MUX2X1 U11891 ( .B(n10347), .A(n10348), .S(N21), .Y(n10346) );
  MUX2X1 U11892 ( .B(n10350), .A(n10351), .S(n10679), .Y(n10349) );
  MUX2X1 U11893 ( .B(n10353), .A(n10354), .S(n10679), .Y(n10352) );
  MUX2X1 U11894 ( .B(n10356), .A(n10357), .S(n10679), .Y(n10355) );
  MUX2X1 U11895 ( .B(n10359), .A(n10360), .S(n10679), .Y(n10358) );
  MUX2X1 U11896 ( .B(n10362), .A(n10363), .S(N21), .Y(n10361) );
  MUX2X1 U11897 ( .B(n10365), .A(n10366), .S(n10680), .Y(n10364) );
  MUX2X1 U11898 ( .B(n10368), .A(n10369), .S(n10680), .Y(n10367) );
  MUX2X1 U11899 ( .B(n10371), .A(n10372), .S(n10680), .Y(n10370) );
  MUX2X1 U11900 ( .B(n10374), .A(n10375), .S(n10680), .Y(n10373) );
  MUX2X1 U11901 ( .B(n10377), .A(n10378), .S(N21), .Y(n10376) );
  MUX2X1 U11902 ( .B(n10380), .A(n10381), .S(n10680), .Y(n10379) );
  MUX2X1 U11903 ( .B(n10383), .A(n10384), .S(n10680), .Y(n10382) );
  MUX2X1 U11904 ( .B(n10386), .A(n10387), .S(n10680), .Y(n10385) );
  MUX2X1 U11905 ( .B(n10389), .A(n10390), .S(n10680), .Y(n10388) );
  MUX2X1 U11906 ( .B(n10392), .A(n10393), .S(N21), .Y(n10391) );
  MUX2X1 U11907 ( .B(n10395), .A(n10396), .S(n10680), .Y(n10394) );
  MUX2X1 U11908 ( .B(n10398), .A(n10399), .S(n10680), .Y(n10397) );
  MUX2X1 U11909 ( .B(n10401), .A(n10402), .S(n10680), .Y(n10400) );
  MUX2X1 U11910 ( .B(n10404), .A(n10405), .S(n10680), .Y(n10403) );
  MUX2X1 U11911 ( .B(n10407), .A(n10408), .S(N21), .Y(n10406) );
  MUX2X1 U11912 ( .B(n10410), .A(n10411), .S(n10681), .Y(n10409) );
  MUX2X1 U11913 ( .B(n10413), .A(n10414), .S(n10681), .Y(n10412) );
  MUX2X1 U11914 ( .B(n10416), .A(n10417), .S(n10681), .Y(n10415) );
  MUX2X1 U11915 ( .B(n10419), .A(n10420), .S(n10681), .Y(n10418) );
  MUX2X1 U11916 ( .B(n10422), .A(n10423), .S(N21), .Y(n10421) );
  MUX2X1 U11917 ( .B(n10425), .A(n10426), .S(n10681), .Y(n10424) );
  MUX2X1 U11918 ( .B(n10428), .A(n10429), .S(n10681), .Y(n10427) );
  MUX2X1 U11919 ( .B(n10431), .A(n10432), .S(n10681), .Y(n10430) );
  MUX2X1 U11920 ( .B(n10434), .A(n10435), .S(n10681), .Y(n10433) );
  MUX2X1 U11921 ( .B(n10437), .A(n10438), .S(N21), .Y(n10436) );
  MUX2X1 U11922 ( .B(n10440), .A(n10441), .S(n10681), .Y(n10439) );
  MUX2X1 U11923 ( .B(n10443), .A(n10444), .S(n10681), .Y(n10442) );
  MUX2X1 U11924 ( .B(n10446), .A(n10447), .S(n10681), .Y(n10445) );
  MUX2X1 U11925 ( .B(n10449), .A(n10450), .S(n10681), .Y(n10448) );
  MUX2X1 U11926 ( .B(n10452), .A(n10453), .S(N21), .Y(n10451) );
  MUX2X1 U11927 ( .B(\RF[30][0] ), .A(\RF[31][0] ), .S(n10538), .Y(n8536) );
  MUX2X1 U11928 ( .B(\RF[28][0] ), .A(\RF[29][0] ), .S(n10538), .Y(n8535) );
  MUX2X1 U11929 ( .B(\RF[26][0] ), .A(\RF[27][0] ), .S(n10538), .Y(n8539) );
  MUX2X1 U11930 ( .B(\RF[24][0] ), .A(\RF[25][0] ), .S(n10538), .Y(n8538) );
  MUX2X1 U11931 ( .B(n8537), .A(n8534), .S(N20), .Y(n8548) );
  MUX2X1 U11932 ( .B(\RF[22][0] ), .A(\RF[23][0] ), .S(n10539), .Y(n8542) );
  MUX2X1 U11933 ( .B(\RF[20][0] ), .A(\RF[21][0] ), .S(n10539), .Y(n8541) );
  MUX2X1 U11934 ( .B(\RF[18][0] ), .A(\RF[19][0] ), .S(n10539), .Y(n8545) );
  MUX2X1 U11935 ( .B(\RF[16][0] ), .A(\RF[17][0] ), .S(n10539), .Y(n8544) );
  MUX2X1 U11936 ( .B(n8543), .A(n8540), .S(N20), .Y(n8547) );
  MUX2X1 U11937 ( .B(\RF[14][0] ), .A(\RF[15][0] ), .S(n10539), .Y(n8551) );
  MUX2X1 U11938 ( .B(\RF[12][0] ), .A(\RF[13][0] ), .S(n10539), .Y(n8550) );
  MUX2X1 U11939 ( .B(\RF[10][0] ), .A(\RF[11][0] ), .S(n10539), .Y(n8554) );
  MUX2X1 U11940 ( .B(\RF[8][0] ), .A(\RF[9][0] ), .S(n10539), .Y(n8553) );
  MUX2X1 U11941 ( .B(n8552), .A(n8549), .S(N20), .Y(n8563) );
  MUX2X1 U11942 ( .B(\RF[6][0] ), .A(\RF[7][0] ), .S(n10539), .Y(n8557) );
  MUX2X1 U11943 ( .B(\RF[4][0] ), .A(\RF[5][0] ), .S(n10539), .Y(n8556) );
  MUX2X1 U11944 ( .B(\RF[2][0] ), .A(\RF[3][0] ), .S(n10539), .Y(n8560) );
  MUX2X1 U11945 ( .B(\RF[0][0] ), .A(\RF[1][0] ), .S(n10539), .Y(n8559) );
  MUX2X1 U11946 ( .B(n8558), .A(n8555), .S(N20), .Y(n8562) );
  MUX2X1 U11947 ( .B(n8561), .A(n8546), .S(N22), .Y(n10454) );
  MUX2X1 U11948 ( .B(\RF[30][1] ), .A(\RF[31][1] ), .S(n10540), .Y(n8566) );
  MUX2X1 U11949 ( .B(\RF[28][1] ), .A(\RF[29][1] ), .S(n10540), .Y(n8565) );
  MUX2X1 U11950 ( .B(\RF[26][1] ), .A(\RF[27][1] ), .S(n10540), .Y(n8569) );
  MUX2X1 U11951 ( .B(\RF[24][1] ), .A(\RF[25][1] ), .S(n10540), .Y(n8568) );
  MUX2X1 U11952 ( .B(n8567), .A(n8564), .S(n10684), .Y(n8578) );
  MUX2X1 U11953 ( .B(\RF[22][1] ), .A(\RF[23][1] ), .S(n10540), .Y(n8572) );
  MUX2X1 U11954 ( .B(\RF[20][1] ), .A(\RF[21][1] ), .S(n10540), .Y(n8571) );
  MUX2X1 U11955 ( .B(\RF[18][1] ), .A(\RF[19][1] ), .S(n10540), .Y(n8575) );
  MUX2X1 U11956 ( .B(\RF[16][1] ), .A(\RF[17][1] ), .S(n10540), .Y(n8574) );
  MUX2X1 U11957 ( .B(n8573), .A(n8570), .S(n10684), .Y(n8577) );
  MUX2X1 U11958 ( .B(\RF[14][1] ), .A(\RF[15][1] ), .S(n10540), .Y(n8581) );
  MUX2X1 U11959 ( .B(\RF[12][1] ), .A(\RF[13][1] ), .S(n10540), .Y(n8580) );
  MUX2X1 U11960 ( .B(\RF[10][1] ), .A(\RF[11][1] ), .S(n10540), .Y(n8584) );
  MUX2X1 U11961 ( .B(\RF[8][1] ), .A(\RF[9][1] ), .S(n10540), .Y(n8583) );
  MUX2X1 U11962 ( .B(n8582), .A(n8579), .S(n10684), .Y(n8593) );
  MUX2X1 U11963 ( .B(\RF[6][1] ), .A(\RF[7][1] ), .S(n10541), .Y(n8587) );
  MUX2X1 U11964 ( .B(\RF[4][1] ), .A(\RF[5][1] ), .S(n10541), .Y(n8586) );
  MUX2X1 U11965 ( .B(\RF[2][1] ), .A(\RF[3][1] ), .S(n10541), .Y(n8590) );
  MUX2X1 U11966 ( .B(\RF[0][1] ), .A(\RF[1][1] ), .S(n10541), .Y(n8589) );
  MUX2X1 U11967 ( .B(n8588), .A(n8585), .S(n10684), .Y(n8592) );
  MUX2X1 U11968 ( .B(n8591), .A(n8576), .S(N22), .Y(n10455) );
  MUX2X1 U11969 ( .B(\RF[30][2] ), .A(\RF[31][2] ), .S(n10541), .Y(n8596) );
  MUX2X1 U11970 ( .B(\RF[28][2] ), .A(\RF[29][2] ), .S(n10541), .Y(n8595) );
  MUX2X1 U11971 ( .B(\RF[26][2] ), .A(\RF[27][2] ), .S(n10541), .Y(n8599) );
  MUX2X1 U11972 ( .B(\RF[24][2] ), .A(\RF[25][2] ), .S(n10541), .Y(n8598) );
  MUX2X1 U11973 ( .B(n8597), .A(n8594), .S(n10684), .Y(n8608) );
  MUX2X1 U11974 ( .B(\RF[22][2] ), .A(\RF[23][2] ), .S(n10541), .Y(n8602) );
  MUX2X1 U11975 ( .B(\RF[20][2] ), .A(\RF[21][2] ), .S(n10541), .Y(n8601) );
  MUX2X1 U11976 ( .B(\RF[18][2] ), .A(\RF[19][2] ), .S(n10541), .Y(n8605) );
  MUX2X1 U11977 ( .B(\RF[16][2] ), .A(\RF[17][2] ), .S(n10541), .Y(n8604) );
  MUX2X1 U11978 ( .B(n8603), .A(n8600), .S(n10684), .Y(n8607) );
  MUX2X1 U11979 ( .B(\RF[14][2] ), .A(\RF[15][2] ), .S(n10542), .Y(n8611) );
  MUX2X1 U11980 ( .B(\RF[12][2] ), .A(\RF[13][2] ), .S(n10542), .Y(n8610) );
  MUX2X1 U11981 ( .B(\RF[10][2] ), .A(\RF[11][2] ), .S(n10542), .Y(n8614) );
  MUX2X1 U11982 ( .B(\RF[8][2] ), .A(\RF[9][2] ), .S(n10542), .Y(n8613) );
  MUX2X1 U11983 ( .B(n8612), .A(n8609), .S(n10684), .Y(n8623) );
  MUX2X1 U11984 ( .B(\RF[6][2] ), .A(\RF[7][2] ), .S(n10542), .Y(n8617) );
  MUX2X1 U11985 ( .B(\RF[4][2] ), .A(\RF[5][2] ), .S(n10542), .Y(n8616) );
  MUX2X1 U11986 ( .B(\RF[2][2] ), .A(\RF[3][2] ), .S(n10542), .Y(n8620) );
  MUX2X1 U11987 ( .B(\RF[0][2] ), .A(\RF[1][2] ), .S(n10542), .Y(n8619) );
  MUX2X1 U11988 ( .B(n8618), .A(n8615), .S(n10684), .Y(n8622) );
  MUX2X1 U11989 ( .B(n8621), .A(n8606), .S(N22), .Y(n10456) );
  MUX2X1 U11990 ( .B(\RF[30][3] ), .A(\RF[31][3] ), .S(n10542), .Y(n8626) );
  MUX2X1 U11991 ( .B(\RF[28][3] ), .A(\RF[29][3] ), .S(n10542), .Y(n8625) );
  MUX2X1 U11992 ( .B(\RF[26][3] ), .A(\RF[27][3] ), .S(n10542), .Y(n8629) );
  MUX2X1 U11993 ( .B(\RF[24][3] ), .A(\RF[25][3] ), .S(n10542), .Y(n8628) );
  MUX2X1 U11994 ( .B(n8627), .A(n8624), .S(n10684), .Y(n8638) );
  MUX2X1 U11995 ( .B(\RF[22][3] ), .A(\RF[23][3] ), .S(n10543), .Y(n8632) );
  MUX2X1 U11996 ( .B(\RF[20][3] ), .A(\RF[21][3] ), .S(n10543), .Y(n8631) );
  MUX2X1 U11997 ( .B(\RF[18][3] ), .A(\RF[19][3] ), .S(n10543), .Y(n8635) );
  MUX2X1 U11998 ( .B(\RF[16][3] ), .A(\RF[17][3] ), .S(n10543), .Y(n8634) );
  MUX2X1 U11999 ( .B(n8633), .A(n8630), .S(n10684), .Y(n8637) );
  MUX2X1 U12000 ( .B(\RF[14][3] ), .A(\RF[15][3] ), .S(n10543), .Y(n8641) );
  MUX2X1 U12001 ( .B(\RF[12][3] ), .A(\RF[13][3] ), .S(n10543), .Y(n8640) );
  MUX2X1 U12002 ( .B(\RF[10][3] ), .A(\RF[11][3] ), .S(n10543), .Y(n8644) );
  MUX2X1 U12003 ( .B(\RF[8][3] ), .A(\RF[9][3] ), .S(n10543), .Y(n8643) );
  MUX2X1 U12004 ( .B(n8642), .A(n8639), .S(n10684), .Y(n8653) );
  MUX2X1 U12005 ( .B(\RF[6][3] ), .A(\RF[7][3] ), .S(n10543), .Y(n8647) );
  MUX2X1 U12006 ( .B(\RF[4][3] ), .A(\RF[5][3] ), .S(n10543), .Y(n8646) );
  MUX2X1 U12007 ( .B(\RF[2][3] ), .A(\RF[3][3] ), .S(n10543), .Y(n8650) );
  MUX2X1 U12008 ( .B(\RF[0][3] ), .A(\RF[1][3] ), .S(n10543), .Y(n8649) );
  MUX2X1 U12009 ( .B(n8648), .A(n8645), .S(n10684), .Y(n8652) );
  MUX2X1 U12010 ( .B(n8651), .A(n8636), .S(N22), .Y(n10457) );
  MUX2X1 U12011 ( .B(\RF[30][4] ), .A(\RF[31][4] ), .S(n10544), .Y(n8656) );
  MUX2X1 U12012 ( .B(\RF[28][4] ), .A(\RF[29][4] ), .S(n10544), .Y(n8655) );
  MUX2X1 U12013 ( .B(\RF[26][4] ), .A(\RF[27][4] ), .S(n10544), .Y(n8659) );
  MUX2X1 U12014 ( .B(\RF[24][4] ), .A(\RF[25][4] ), .S(n10544), .Y(n8658) );
  MUX2X1 U12015 ( .B(n8657), .A(n8654), .S(n10685), .Y(n8668) );
  MUX2X1 U12016 ( .B(\RF[22][4] ), .A(\RF[23][4] ), .S(n10544), .Y(n8662) );
  MUX2X1 U12017 ( .B(\RF[20][4] ), .A(\RF[21][4] ), .S(n10544), .Y(n8661) );
  MUX2X1 U12018 ( .B(\RF[18][4] ), .A(\RF[19][4] ), .S(n10544), .Y(n8665) );
  MUX2X1 U12019 ( .B(\RF[16][4] ), .A(\RF[17][4] ), .S(n10544), .Y(n8664) );
  MUX2X1 U12020 ( .B(n8663), .A(n8660), .S(n10685), .Y(n8667) );
  MUX2X1 U12021 ( .B(\RF[14][4] ), .A(\RF[15][4] ), .S(n10544), .Y(n8671) );
  MUX2X1 U12022 ( .B(\RF[12][4] ), .A(\RF[13][4] ), .S(n10544), .Y(n8670) );
  MUX2X1 U12023 ( .B(\RF[10][4] ), .A(\RF[11][4] ), .S(n10544), .Y(n8674) );
  MUX2X1 U12024 ( .B(\RF[8][4] ), .A(\RF[9][4] ), .S(n10544), .Y(n8673) );
  MUX2X1 U12025 ( .B(n8672), .A(n8669), .S(n10685), .Y(n8683) );
  MUX2X1 U12026 ( .B(\RF[6][4] ), .A(\RF[7][4] ), .S(n10545), .Y(n8677) );
  MUX2X1 U12027 ( .B(\RF[4][4] ), .A(\RF[5][4] ), .S(n10545), .Y(n8676) );
  MUX2X1 U12028 ( .B(\RF[2][4] ), .A(\RF[3][4] ), .S(n10545), .Y(n8680) );
  MUX2X1 U12029 ( .B(\RF[0][4] ), .A(\RF[1][4] ), .S(n10545), .Y(n8679) );
  MUX2X1 U12030 ( .B(n8678), .A(n8675), .S(n10685), .Y(n8682) );
  MUX2X1 U12031 ( .B(n8681), .A(n8666), .S(N22), .Y(n10458) );
  MUX2X1 U12032 ( .B(\RF[30][5] ), .A(\RF[31][5] ), .S(n10545), .Y(n8686) );
  MUX2X1 U12033 ( .B(\RF[28][5] ), .A(\RF[29][5] ), .S(n10545), .Y(n8685) );
  MUX2X1 U12034 ( .B(\RF[26][5] ), .A(\RF[27][5] ), .S(n10545), .Y(n8689) );
  MUX2X1 U12035 ( .B(\RF[24][5] ), .A(\RF[25][5] ), .S(n10545), .Y(n8688) );
  MUX2X1 U12036 ( .B(n8687), .A(n8684), .S(n10685), .Y(n8698) );
  MUX2X1 U12037 ( .B(\RF[22][5] ), .A(\RF[23][5] ), .S(n10545), .Y(n8692) );
  MUX2X1 U12038 ( .B(\RF[20][5] ), .A(\RF[21][5] ), .S(n10545), .Y(n8691) );
  MUX2X1 U12039 ( .B(\RF[18][5] ), .A(\RF[19][5] ), .S(n10545), .Y(n8695) );
  MUX2X1 U12040 ( .B(\RF[16][5] ), .A(\RF[17][5] ), .S(n10545), .Y(n8694) );
  MUX2X1 U12041 ( .B(n8693), .A(n8690), .S(n10685), .Y(n8697) );
  MUX2X1 U12042 ( .B(\RF[14][5] ), .A(\RF[15][5] ), .S(n10546), .Y(n8701) );
  MUX2X1 U12043 ( .B(\RF[12][5] ), .A(\RF[13][5] ), .S(n10546), .Y(n8700) );
  MUX2X1 U12044 ( .B(\RF[10][5] ), .A(\RF[11][5] ), .S(n10546), .Y(n8704) );
  MUX2X1 U12045 ( .B(\RF[8][5] ), .A(\RF[9][5] ), .S(n10546), .Y(n8703) );
  MUX2X1 U12046 ( .B(n8702), .A(n8699), .S(n10685), .Y(n8713) );
  MUX2X1 U12047 ( .B(\RF[6][5] ), .A(\RF[7][5] ), .S(n10546), .Y(n8707) );
  MUX2X1 U12048 ( .B(\RF[4][5] ), .A(\RF[5][5] ), .S(n10546), .Y(n8706) );
  MUX2X1 U12049 ( .B(\RF[2][5] ), .A(\RF[3][5] ), .S(n10546), .Y(n8710) );
  MUX2X1 U12050 ( .B(\RF[0][5] ), .A(\RF[1][5] ), .S(n10546), .Y(n8709) );
  MUX2X1 U12051 ( .B(n8708), .A(n8705), .S(n10685), .Y(n8712) );
  MUX2X1 U12052 ( .B(n8711), .A(n8696), .S(N22), .Y(n10459) );
  MUX2X1 U12053 ( .B(\RF[30][6] ), .A(\RF[31][6] ), .S(n10546), .Y(n8716) );
  MUX2X1 U12054 ( .B(\RF[28][6] ), .A(\RF[29][6] ), .S(n10546), .Y(n8715) );
  MUX2X1 U12055 ( .B(\RF[26][6] ), .A(\RF[27][6] ), .S(n10546), .Y(n8719) );
  MUX2X1 U12056 ( .B(\RF[24][6] ), .A(\RF[25][6] ), .S(n10546), .Y(n8718) );
  MUX2X1 U12057 ( .B(n8717), .A(n8714), .S(n10685), .Y(n8728) );
  MUX2X1 U12058 ( .B(\RF[22][6] ), .A(\RF[23][6] ), .S(n10547), .Y(n8722) );
  MUX2X1 U12059 ( .B(\RF[20][6] ), .A(\RF[21][6] ), .S(n10547), .Y(n8721) );
  MUX2X1 U12060 ( .B(\RF[18][6] ), .A(\RF[19][6] ), .S(n10547), .Y(n8725) );
  MUX2X1 U12061 ( .B(\RF[16][6] ), .A(\RF[17][6] ), .S(n10547), .Y(n8724) );
  MUX2X1 U12062 ( .B(n8723), .A(n8720), .S(n10685), .Y(n8727) );
  MUX2X1 U12063 ( .B(\RF[14][6] ), .A(\RF[15][6] ), .S(n10547), .Y(n8731) );
  MUX2X1 U12064 ( .B(\RF[12][6] ), .A(\RF[13][6] ), .S(n10547), .Y(n8730) );
  MUX2X1 U12065 ( .B(\RF[10][6] ), .A(\RF[11][6] ), .S(n10547), .Y(n8734) );
  MUX2X1 U12066 ( .B(\RF[8][6] ), .A(\RF[9][6] ), .S(n10547), .Y(n8733) );
  MUX2X1 U12067 ( .B(n8732), .A(n8729), .S(n10685), .Y(n8743) );
  MUX2X1 U12068 ( .B(\RF[6][6] ), .A(\RF[7][6] ), .S(n10547), .Y(n8737) );
  MUX2X1 U12069 ( .B(\RF[4][6] ), .A(\RF[5][6] ), .S(n10547), .Y(n8736) );
  MUX2X1 U12070 ( .B(\RF[2][6] ), .A(\RF[3][6] ), .S(n10547), .Y(n8740) );
  MUX2X1 U12071 ( .B(\RF[0][6] ), .A(\RF[1][6] ), .S(n10547), .Y(n8739) );
  MUX2X1 U12072 ( .B(n8738), .A(n8735), .S(n10685), .Y(n8742) );
  MUX2X1 U12073 ( .B(n8741), .A(n8726), .S(N22), .Y(n10460) );
  MUX2X1 U12074 ( .B(\RF[30][7] ), .A(\RF[31][7] ), .S(n10548), .Y(n8746) );
  MUX2X1 U12075 ( .B(\RF[28][7] ), .A(\RF[29][7] ), .S(n10548), .Y(n8745) );
  MUX2X1 U12076 ( .B(\RF[26][7] ), .A(\RF[27][7] ), .S(n10548), .Y(n8749) );
  MUX2X1 U12077 ( .B(\RF[24][7] ), .A(\RF[25][7] ), .S(n10548), .Y(n8748) );
  MUX2X1 U12078 ( .B(n8747), .A(n8744), .S(n10686), .Y(n8758) );
  MUX2X1 U12079 ( .B(\RF[22][7] ), .A(\RF[23][7] ), .S(n10548), .Y(n8752) );
  MUX2X1 U12080 ( .B(\RF[20][7] ), .A(\RF[21][7] ), .S(n10548), .Y(n8751) );
  MUX2X1 U12081 ( .B(\RF[18][7] ), .A(\RF[19][7] ), .S(n10548), .Y(n8755) );
  MUX2X1 U12082 ( .B(\RF[16][7] ), .A(\RF[17][7] ), .S(n10548), .Y(n8754) );
  MUX2X1 U12083 ( .B(n8753), .A(n8750), .S(n10686), .Y(n8757) );
  MUX2X1 U12084 ( .B(\RF[14][7] ), .A(\RF[15][7] ), .S(n10548), .Y(n8761) );
  MUX2X1 U12085 ( .B(\RF[12][7] ), .A(\RF[13][7] ), .S(n10548), .Y(n8760) );
  MUX2X1 U12086 ( .B(\RF[10][7] ), .A(\RF[11][7] ), .S(n10548), .Y(n8764) );
  MUX2X1 U12087 ( .B(\RF[8][7] ), .A(\RF[9][7] ), .S(n10548), .Y(n8763) );
  MUX2X1 U12088 ( .B(n8762), .A(n8759), .S(n10686), .Y(n8773) );
  MUX2X1 U12089 ( .B(\RF[6][7] ), .A(\RF[7][7] ), .S(n10549), .Y(n8767) );
  MUX2X1 U12090 ( .B(\RF[4][7] ), .A(\RF[5][7] ), .S(n10549), .Y(n8766) );
  MUX2X1 U12091 ( .B(\RF[2][7] ), .A(\RF[3][7] ), .S(n10549), .Y(n8770) );
  MUX2X1 U12092 ( .B(\RF[0][7] ), .A(\RF[1][7] ), .S(n10549), .Y(n8769) );
  MUX2X1 U12093 ( .B(n8768), .A(n8765), .S(n10686), .Y(n8772) );
  MUX2X1 U12094 ( .B(n8771), .A(n8756), .S(N22), .Y(n10461) );
  MUX2X1 U12095 ( .B(\RF[30][8] ), .A(\RF[31][8] ), .S(n10549), .Y(n8776) );
  MUX2X1 U12096 ( .B(\RF[28][8] ), .A(\RF[29][8] ), .S(n10549), .Y(n8775) );
  MUX2X1 U12097 ( .B(\RF[26][8] ), .A(\RF[27][8] ), .S(n10549), .Y(n8779) );
  MUX2X1 U12098 ( .B(\RF[24][8] ), .A(\RF[25][8] ), .S(n10549), .Y(n8778) );
  MUX2X1 U12099 ( .B(n8777), .A(n8774), .S(n10686), .Y(n8788) );
  MUX2X1 U12100 ( .B(\RF[22][8] ), .A(\RF[23][8] ), .S(n10549), .Y(n8782) );
  MUX2X1 U12101 ( .B(\RF[20][8] ), .A(\RF[21][8] ), .S(n10549), .Y(n8781) );
  MUX2X1 U12102 ( .B(\RF[18][8] ), .A(\RF[19][8] ), .S(n10549), .Y(n8785) );
  MUX2X1 U12103 ( .B(\RF[16][8] ), .A(\RF[17][8] ), .S(n10549), .Y(n8784) );
  MUX2X1 U12104 ( .B(n8783), .A(n8780), .S(n10686), .Y(n8787) );
  MUX2X1 U12105 ( .B(\RF[14][8] ), .A(\RF[15][8] ), .S(n10550), .Y(n8791) );
  MUX2X1 U12106 ( .B(\RF[12][8] ), .A(\RF[13][8] ), .S(n10550), .Y(n8790) );
  MUX2X1 U12107 ( .B(\RF[10][8] ), .A(\RF[11][8] ), .S(n10550), .Y(n8794) );
  MUX2X1 U12108 ( .B(\RF[8][8] ), .A(\RF[9][8] ), .S(n10550), .Y(n8793) );
  MUX2X1 U12109 ( .B(n8792), .A(n8789), .S(n10686), .Y(n8803) );
  MUX2X1 U12110 ( .B(\RF[6][8] ), .A(\RF[7][8] ), .S(n10550), .Y(n8797) );
  MUX2X1 U12111 ( .B(\RF[4][8] ), .A(\RF[5][8] ), .S(n10550), .Y(n8796) );
  MUX2X1 U12112 ( .B(\RF[2][8] ), .A(\RF[3][8] ), .S(n10550), .Y(n8800) );
  MUX2X1 U12113 ( .B(\RF[0][8] ), .A(\RF[1][8] ), .S(n10550), .Y(n8799) );
  MUX2X1 U12114 ( .B(n8798), .A(n8795), .S(n10686), .Y(n8802) );
  MUX2X1 U12115 ( .B(n8801), .A(n8786), .S(N22), .Y(n10462) );
  MUX2X1 U12116 ( .B(\RF[30][9] ), .A(\RF[31][9] ), .S(n10550), .Y(n8806) );
  MUX2X1 U12117 ( .B(\RF[28][9] ), .A(\RF[29][9] ), .S(n10550), .Y(n8805) );
  MUX2X1 U12118 ( .B(\RF[26][9] ), .A(\RF[27][9] ), .S(n10550), .Y(n8809) );
  MUX2X1 U12119 ( .B(\RF[24][9] ), .A(\RF[25][9] ), .S(n10550), .Y(n8808) );
  MUX2X1 U12120 ( .B(n8807), .A(n8804), .S(n10686), .Y(n8818) );
  MUX2X1 U12121 ( .B(\RF[22][9] ), .A(\RF[23][9] ), .S(n10551), .Y(n8812) );
  MUX2X1 U12122 ( .B(\RF[20][9] ), .A(\RF[21][9] ), .S(n10551), .Y(n8811) );
  MUX2X1 U12123 ( .B(\RF[18][9] ), .A(\RF[19][9] ), .S(n10551), .Y(n8815) );
  MUX2X1 U12124 ( .B(\RF[16][9] ), .A(\RF[17][9] ), .S(n10551), .Y(n8814) );
  MUX2X1 U12125 ( .B(n8813), .A(n8810), .S(n10686), .Y(n8817) );
  MUX2X1 U12126 ( .B(\RF[14][9] ), .A(\RF[15][9] ), .S(n10551), .Y(n8821) );
  MUX2X1 U12127 ( .B(\RF[12][9] ), .A(\RF[13][9] ), .S(n10551), .Y(n8820) );
  MUX2X1 U12128 ( .B(\RF[10][9] ), .A(\RF[11][9] ), .S(n10551), .Y(n8824) );
  MUX2X1 U12129 ( .B(\RF[8][9] ), .A(\RF[9][9] ), .S(n10551), .Y(n8823) );
  MUX2X1 U12130 ( .B(n8822), .A(n8819), .S(n10686), .Y(n8833) );
  MUX2X1 U12131 ( .B(\RF[6][9] ), .A(\RF[7][9] ), .S(n10551), .Y(n8827) );
  MUX2X1 U12132 ( .B(\RF[4][9] ), .A(\RF[5][9] ), .S(n10551), .Y(n8826) );
  MUX2X1 U12133 ( .B(\RF[2][9] ), .A(\RF[3][9] ), .S(n10551), .Y(n8830) );
  MUX2X1 U12134 ( .B(\RF[0][9] ), .A(\RF[1][9] ), .S(n10551), .Y(n8829) );
  MUX2X1 U12135 ( .B(n8828), .A(n8825), .S(n10686), .Y(n8832) );
  MUX2X1 U12136 ( .B(n8831), .A(n8816), .S(N22), .Y(n10463) );
  MUX2X1 U12137 ( .B(\RF[30][10] ), .A(\RF[31][10] ), .S(n10552), .Y(n8836) );
  MUX2X1 U12138 ( .B(\RF[28][10] ), .A(\RF[29][10] ), .S(n10552), .Y(n8835) );
  MUX2X1 U12139 ( .B(\RF[26][10] ), .A(\RF[27][10] ), .S(n10552), .Y(n8839) );
  MUX2X1 U12140 ( .B(\RF[24][10] ), .A(\RF[25][10] ), .S(n10552), .Y(n8838) );
  MUX2X1 U12141 ( .B(n8837), .A(n8834), .S(n10687), .Y(n8848) );
  MUX2X1 U12142 ( .B(\RF[22][10] ), .A(\RF[23][10] ), .S(n10552), .Y(n8842) );
  MUX2X1 U12143 ( .B(\RF[20][10] ), .A(\RF[21][10] ), .S(n10552), .Y(n8841) );
  MUX2X1 U12144 ( .B(\RF[18][10] ), .A(\RF[19][10] ), .S(n10552), .Y(n8845) );
  MUX2X1 U12145 ( .B(\RF[16][10] ), .A(\RF[17][10] ), .S(n10552), .Y(n8844) );
  MUX2X1 U12146 ( .B(n8843), .A(n8840), .S(n10687), .Y(n8847) );
  MUX2X1 U12147 ( .B(\RF[14][10] ), .A(\RF[15][10] ), .S(n10552), .Y(n8851) );
  MUX2X1 U12148 ( .B(\RF[12][10] ), .A(\RF[13][10] ), .S(n10552), .Y(n8850) );
  MUX2X1 U12149 ( .B(\RF[10][10] ), .A(\RF[11][10] ), .S(n10552), .Y(n8854) );
  MUX2X1 U12150 ( .B(\RF[8][10] ), .A(\RF[9][10] ), .S(n10552), .Y(n8853) );
  MUX2X1 U12151 ( .B(n8852), .A(n8849), .S(n10687), .Y(n8863) );
  MUX2X1 U12152 ( .B(\RF[6][10] ), .A(\RF[7][10] ), .S(n10553), .Y(n8857) );
  MUX2X1 U12153 ( .B(\RF[4][10] ), .A(\RF[5][10] ), .S(n10553), .Y(n8856) );
  MUX2X1 U12154 ( .B(\RF[2][10] ), .A(\RF[3][10] ), .S(n10553), .Y(n8860) );
  MUX2X1 U12155 ( .B(\RF[0][10] ), .A(\RF[1][10] ), .S(n10553), .Y(n8859) );
  MUX2X1 U12156 ( .B(n8858), .A(n8855), .S(n10687), .Y(n8862) );
  MUX2X1 U12157 ( .B(n8861), .A(n8846), .S(N22), .Y(n10464) );
  MUX2X1 U12158 ( .B(\RF[30][11] ), .A(\RF[31][11] ), .S(n10553), .Y(n8866) );
  MUX2X1 U12159 ( .B(\RF[28][11] ), .A(\RF[29][11] ), .S(n10553), .Y(n8865) );
  MUX2X1 U12160 ( .B(\RF[26][11] ), .A(\RF[27][11] ), .S(n10553), .Y(n8869) );
  MUX2X1 U12161 ( .B(\RF[24][11] ), .A(\RF[25][11] ), .S(n10553), .Y(n8868) );
  MUX2X1 U12162 ( .B(n8867), .A(n8864), .S(n10687), .Y(n8878) );
  MUX2X1 U12163 ( .B(\RF[22][11] ), .A(\RF[23][11] ), .S(n10553), .Y(n8872) );
  MUX2X1 U12164 ( .B(\RF[20][11] ), .A(\RF[21][11] ), .S(n10553), .Y(n8871) );
  MUX2X1 U12165 ( .B(\RF[18][11] ), .A(\RF[19][11] ), .S(n10553), .Y(n8875) );
  MUX2X1 U12166 ( .B(\RF[16][11] ), .A(\RF[17][11] ), .S(n10553), .Y(n8874) );
  MUX2X1 U12167 ( .B(n8873), .A(n8870), .S(n10687), .Y(n8877) );
  MUX2X1 U12168 ( .B(\RF[14][11] ), .A(\RF[15][11] ), .S(n10554), .Y(n8881) );
  MUX2X1 U12169 ( .B(\RF[12][11] ), .A(\RF[13][11] ), .S(n10554), .Y(n8880) );
  MUX2X1 U12170 ( .B(\RF[10][11] ), .A(\RF[11][11] ), .S(n10554), .Y(n8884) );
  MUX2X1 U12171 ( .B(\RF[8][11] ), .A(\RF[9][11] ), .S(n10554), .Y(n8883) );
  MUX2X1 U12172 ( .B(n8882), .A(n8879), .S(n10687), .Y(n8893) );
  MUX2X1 U12173 ( .B(\RF[6][11] ), .A(\RF[7][11] ), .S(n10554), .Y(n8887) );
  MUX2X1 U12174 ( .B(\RF[4][11] ), .A(\RF[5][11] ), .S(n10554), .Y(n8886) );
  MUX2X1 U12175 ( .B(\RF[2][11] ), .A(\RF[3][11] ), .S(n10554), .Y(n8890) );
  MUX2X1 U12176 ( .B(\RF[0][11] ), .A(\RF[1][11] ), .S(n10554), .Y(n8889) );
  MUX2X1 U12177 ( .B(n8888), .A(n8885), .S(n10687), .Y(n8892) );
  MUX2X1 U12178 ( .B(n8891), .A(n8876), .S(N22), .Y(n10465) );
  MUX2X1 U12179 ( .B(\RF[30][12] ), .A(\RF[31][12] ), .S(n10554), .Y(n8896) );
  MUX2X1 U12180 ( .B(\RF[28][12] ), .A(\RF[29][12] ), .S(n10554), .Y(n8895) );
  MUX2X1 U12181 ( .B(\RF[26][12] ), .A(\RF[27][12] ), .S(n10554), .Y(n8899) );
  MUX2X1 U12182 ( .B(\RF[24][12] ), .A(\RF[25][12] ), .S(n10554), .Y(n8898) );
  MUX2X1 U12183 ( .B(n8897), .A(n8894), .S(n10687), .Y(n8908) );
  MUX2X1 U12184 ( .B(\RF[22][12] ), .A(\RF[23][12] ), .S(n10555), .Y(n8902) );
  MUX2X1 U12185 ( .B(\RF[20][12] ), .A(\RF[21][12] ), .S(n10555), .Y(n8901) );
  MUX2X1 U12186 ( .B(\RF[18][12] ), .A(\RF[19][12] ), .S(n10555), .Y(n8905) );
  MUX2X1 U12187 ( .B(\RF[16][12] ), .A(\RF[17][12] ), .S(n10555), .Y(n8904) );
  MUX2X1 U12188 ( .B(n8903), .A(n8900), .S(n10687), .Y(n8907) );
  MUX2X1 U12189 ( .B(\RF[14][12] ), .A(\RF[15][12] ), .S(n10555), .Y(n8911) );
  MUX2X1 U12190 ( .B(\RF[12][12] ), .A(\RF[13][12] ), .S(n10555), .Y(n8910) );
  MUX2X1 U12191 ( .B(\RF[10][12] ), .A(\RF[11][12] ), .S(n10555), .Y(n8914) );
  MUX2X1 U12192 ( .B(\RF[8][12] ), .A(\RF[9][12] ), .S(n10555), .Y(n8913) );
  MUX2X1 U12193 ( .B(n8912), .A(n8909), .S(n10687), .Y(n8923) );
  MUX2X1 U12194 ( .B(\RF[6][12] ), .A(\RF[7][12] ), .S(n10555), .Y(n8917) );
  MUX2X1 U12195 ( .B(\RF[4][12] ), .A(\RF[5][12] ), .S(n10555), .Y(n8916) );
  MUX2X1 U12196 ( .B(\RF[2][12] ), .A(\RF[3][12] ), .S(n10555), .Y(n8920) );
  MUX2X1 U12197 ( .B(\RF[0][12] ), .A(\RF[1][12] ), .S(n10555), .Y(n8919) );
  MUX2X1 U12198 ( .B(n8918), .A(n8915), .S(n10687), .Y(n8922) );
  MUX2X1 U12199 ( .B(n8921), .A(n8906), .S(N22), .Y(n10466) );
  MUX2X1 U12200 ( .B(\RF[30][13] ), .A(\RF[31][13] ), .S(n10556), .Y(n8926) );
  MUX2X1 U12201 ( .B(\RF[28][13] ), .A(\RF[29][13] ), .S(n10556), .Y(n8925) );
  MUX2X1 U12202 ( .B(\RF[26][13] ), .A(\RF[27][13] ), .S(n10556), .Y(n8929) );
  MUX2X1 U12203 ( .B(\RF[24][13] ), .A(\RF[25][13] ), .S(n10556), .Y(n8928) );
  MUX2X1 U12204 ( .B(n8927), .A(n8924), .S(n10686), .Y(n8938) );
  MUX2X1 U12205 ( .B(\RF[22][13] ), .A(\RF[23][13] ), .S(n10556), .Y(n8932) );
  MUX2X1 U12206 ( .B(\RF[20][13] ), .A(\RF[21][13] ), .S(n10556), .Y(n8931) );
  MUX2X1 U12207 ( .B(\RF[18][13] ), .A(\RF[19][13] ), .S(n10556), .Y(n8935) );
  MUX2X1 U12208 ( .B(\RF[16][13] ), .A(\RF[17][13] ), .S(n10556), .Y(n8934) );
  MUX2X1 U12209 ( .B(n8933), .A(n8930), .S(n10687), .Y(n8937) );
  MUX2X1 U12210 ( .B(\RF[14][13] ), .A(\RF[15][13] ), .S(n10556), .Y(n8941) );
  MUX2X1 U12211 ( .B(\RF[12][13] ), .A(\RF[13][13] ), .S(n10556), .Y(n8940) );
  MUX2X1 U12212 ( .B(\RF[10][13] ), .A(\RF[11][13] ), .S(n10556), .Y(n8944) );
  MUX2X1 U12213 ( .B(\RF[8][13] ), .A(\RF[9][13] ), .S(n10556), .Y(n8943) );
  MUX2X1 U12214 ( .B(n8942), .A(n8939), .S(N20), .Y(n8953) );
  MUX2X1 U12215 ( .B(\RF[6][13] ), .A(\RF[7][13] ), .S(n10557), .Y(n8947) );
  MUX2X1 U12216 ( .B(\RF[4][13] ), .A(\RF[5][13] ), .S(n10557), .Y(n8946) );
  MUX2X1 U12217 ( .B(\RF[2][13] ), .A(\RF[3][13] ), .S(n10557), .Y(n8950) );
  MUX2X1 U12218 ( .B(\RF[0][13] ), .A(\RF[1][13] ), .S(n10557), .Y(n8949) );
  MUX2X1 U12219 ( .B(n8948), .A(n8945), .S(n10692), .Y(n8952) );
  MUX2X1 U12220 ( .B(n8951), .A(n8936), .S(N22), .Y(n10467) );
  MUX2X1 U12221 ( .B(\RF[30][14] ), .A(\RF[31][14] ), .S(n10557), .Y(n8956) );
  MUX2X1 U12222 ( .B(\RF[28][14] ), .A(\RF[29][14] ), .S(n10557), .Y(n8955) );
  MUX2X1 U12223 ( .B(\RF[26][14] ), .A(\RF[27][14] ), .S(n10557), .Y(n8959) );
  MUX2X1 U12224 ( .B(\RF[24][14] ), .A(\RF[25][14] ), .S(n10557), .Y(n8958) );
  MUX2X1 U12225 ( .B(n8957), .A(n8954), .S(n10697), .Y(n8968) );
  MUX2X1 U12226 ( .B(\RF[22][14] ), .A(\RF[23][14] ), .S(n10557), .Y(n8962) );
  MUX2X1 U12227 ( .B(\RF[20][14] ), .A(\RF[21][14] ), .S(n10557), .Y(n8961) );
  MUX2X1 U12228 ( .B(\RF[18][14] ), .A(\RF[19][14] ), .S(n10557), .Y(n8965) );
  MUX2X1 U12229 ( .B(\RF[16][14] ), .A(\RF[17][14] ), .S(n10557), .Y(n8964) );
  MUX2X1 U12230 ( .B(n8963), .A(n8960), .S(n10689), .Y(n8967) );
  MUX2X1 U12231 ( .B(\RF[14][14] ), .A(\RF[15][14] ), .S(n10558), .Y(n8971) );
  MUX2X1 U12232 ( .B(\RF[12][14] ), .A(\RF[13][14] ), .S(n10558), .Y(n8970) );
  MUX2X1 U12233 ( .B(\RF[10][14] ), .A(\RF[11][14] ), .S(n10558), .Y(n8974) );
  MUX2X1 U12234 ( .B(\RF[8][14] ), .A(\RF[9][14] ), .S(n10558), .Y(n8973) );
  MUX2X1 U12235 ( .B(n8972), .A(n8969), .S(n10698), .Y(n8983) );
  MUX2X1 U12236 ( .B(\RF[6][14] ), .A(\RF[7][14] ), .S(n10558), .Y(n8977) );
  MUX2X1 U12237 ( .B(\RF[4][14] ), .A(\RF[5][14] ), .S(n10558), .Y(n8976) );
  MUX2X1 U12238 ( .B(\RF[2][14] ), .A(\RF[3][14] ), .S(n10558), .Y(n8980) );
  MUX2X1 U12239 ( .B(\RF[0][14] ), .A(\RF[1][14] ), .S(n10558), .Y(n8979) );
  MUX2X1 U12240 ( .B(n8978), .A(n8975), .S(n10693), .Y(n8982) );
  MUX2X1 U12241 ( .B(n8981), .A(n8966), .S(N22), .Y(n10468) );
  MUX2X1 U12242 ( .B(\RF[30][15] ), .A(\RF[31][15] ), .S(n10558), .Y(n8986) );
  MUX2X1 U12243 ( .B(\RF[28][15] ), .A(\RF[29][15] ), .S(n10558), .Y(n8985) );
  MUX2X1 U12244 ( .B(\RF[26][15] ), .A(\RF[27][15] ), .S(n10558), .Y(n8989) );
  MUX2X1 U12245 ( .B(\RF[24][15] ), .A(\RF[25][15] ), .S(n10558), .Y(n8988) );
  MUX2X1 U12246 ( .B(n8987), .A(n8984), .S(n10695), .Y(n8998) );
  MUX2X1 U12247 ( .B(\RF[22][15] ), .A(\RF[23][15] ), .S(n10559), .Y(n8992) );
  MUX2X1 U12248 ( .B(\RF[20][15] ), .A(\RF[21][15] ), .S(n10559), .Y(n8991) );
  MUX2X1 U12249 ( .B(\RF[18][15] ), .A(\RF[19][15] ), .S(n10559), .Y(n8995) );
  MUX2X1 U12250 ( .B(\RF[16][15] ), .A(\RF[17][15] ), .S(n10559), .Y(n8994) );
  MUX2X1 U12251 ( .B(n8993), .A(n8990), .S(n10699), .Y(n8997) );
  MUX2X1 U12252 ( .B(\RF[14][15] ), .A(\RF[15][15] ), .S(n10559), .Y(n9001) );
  MUX2X1 U12253 ( .B(\RF[12][15] ), .A(\RF[13][15] ), .S(n10559), .Y(n9000) );
  MUX2X1 U12254 ( .B(\RF[10][15] ), .A(\RF[11][15] ), .S(n10559), .Y(n9004) );
  MUX2X1 U12255 ( .B(\RF[8][15] ), .A(\RF[9][15] ), .S(n10559), .Y(n9003) );
  MUX2X1 U12256 ( .B(n9002), .A(n8999), .S(n10700), .Y(n9013) );
  MUX2X1 U12257 ( .B(\RF[6][15] ), .A(\RF[7][15] ), .S(n10559), .Y(n9007) );
  MUX2X1 U12258 ( .B(\RF[4][15] ), .A(\RF[5][15] ), .S(n10559), .Y(n9006) );
  MUX2X1 U12259 ( .B(\RF[2][15] ), .A(\RF[3][15] ), .S(n10559), .Y(n9010) );
  MUX2X1 U12260 ( .B(\RF[0][15] ), .A(\RF[1][15] ), .S(n10559), .Y(n9009) );
  MUX2X1 U12261 ( .B(n9008), .A(n9005), .S(n10684), .Y(n9012) );
  MUX2X1 U12262 ( .B(n9011), .A(n8996), .S(N22), .Y(n10469) );
  MUX2X1 U12263 ( .B(\RF[30][16] ), .A(\RF[31][16] ), .S(n10560), .Y(n9016) );
  MUX2X1 U12264 ( .B(\RF[28][16] ), .A(\RF[29][16] ), .S(n10560), .Y(n9015) );
  MUX2X1 U12265 ( .B(\RF[26][16] ), .A(\RF[27][16] ), .S(n10560), .Y(n9019) );
  MUX2X1 U12266 ( .B(\RF[24][16] ), .A(\RF[25][16] ), .S(n10560), .Y(n9018) );
  MUX2X1 U12267 ( .B(n9017), .A(n9014), .S(n10688), .Y(n9028) );
  MUX2X1 U12268 ( .B(\RF[22][16] ), .A(\RF[23][16] ), .S(n10560), .Y(n9022) );
  MUX2X1 U12269 ( .B(\RF[20][16] ), .A(\RF[21][16] ), .S(n10560), .Y(n9021) );
  MUX2X1 U12270 ( .B(\RF[18][16] ), .A(\RF[19][16] ), .S(n10560), .Y(n9025) );
  MUX2X1 U12271 ( .B(\RF[16][16] ), .A(\RF[17][16] ), .S(n10560), .Y(n9024) );
  MUX2X1 U12272 ( .B(n9023), .A(n9020), .S(n10688), .Y(n9027) );
  MUX2X1 U12273 ( .B(\RF[14][16] ), .A(\RF[15][16] ), .S(n10560), .Y(n9031) );
  MUX2X1 U12274 ( .B(\RF[12][16] ), .A(\RF[13][16] ), .S(n10560), .Y(n9030) );
  MUX2X1 U12275 ( .B(\RF[10][16] ), .A(\RF[11][16] ), .S(n10560), .Y(n9034) );
  MUX2X1 U12276 ( .B(\RF[8][16] ), .A(\RF[9][16] ), .S(n10560), .Y(n9033) );
  MUX2X1 U12277 ( .B(n9032), .A(n9029), .S(n10688), .Y(n9043) );
  MUX2X1 U12278 ( .B(\RF[6][16] ), .A(\RF[7][16] ), .S(n10561), .Y(n9037) );
  MUX2X1 U12279 ( .B(\RF[4][16] ), .A(\RF[5][16] ), .S(n10561), .Y(n9036) );
  MUX2X1 U12280 ( .B(\RF[2][16] ), .A(\RF[3][16] ), .S(n10561), .Y(n9040) );
  MUX2X1 U12281 ( .B(\RF[0][16] ), .A(\RF[1][16] ), .S(n10561), .Y(n9039) );
  MUX2X1 U12282 ( .B(n9038), .A(n9035), .S(n10688), .Y(n9042) );
  MUX2X1 U12283 ( .B(n9041), .A(n9026), .S(N22), .Y(n10470) );
  MUX2X1 U12284 ( .B(\RF[30][17] ), .A(\RF[31][17] ), .S(n10561), .Y(n9046) );
  MUX2X1 U12285 ( .B(\RF[28][17] ), .A(\RF[29][17] ), .S(n10561), .Y(n9045) );
  MUX2X1 U12286 ( .B(\RF[26][17] ), .A(\RF[27][17] ), .S(n10561), .Y(n9049) );
  MUX2X1 U12287 ( .B(\RF[24][17] ), .A(\RF[25][17] ), .S(n10561), .Y(n9048) );
  MUX2X1 U12288 ( .B(n9047), .A(n9044), .S(n10688), .Y(n9058) );
  MUX2X1 U12289 ( .B(\RF[22][17] ), .A(\RF[23][17] ), .S(n10561), .Y(n9052) );
  MUX2X1 U12290 ( .B(\RF[20][17] ), .A(\RF[21][17] ), .S(n10561), .Y(n9051) );
  MUX2X1 U12291 ( .B(\RF[18][17] ), .A(\RF[19][17] ), .S(n10561), .Y(n9055) );
  MUX2X1 U12292 ( .B(\RF[16][17] ), .A(\RF[17][17] ), .S(n10561), .Y(n9054) );
  MUX2X1 U12293 ( .B(n9053), .A(n9050), .S(n10688), .Y(n9057) );
  MUX2X1 U12294 ( .B(\RF[14][17] ), .A(\RF[15][17] ), .S(n10562), .Y(n9061) );
  MUX2X1 U12295 ( .B(\RF[12][17] ), .A(\RF[13][17] ), .S(n10562), .Y(n9060) );
  MUX2X1 U12296 ( .B(\RF[10][17] ), .A(\RF[11][17] ), .S(n10562), .Y(n9064) );
  MUX2X1 U12297 ( .B(\RF[8][17] ), .A(\RF[9][17] ), .S(n10562), .Y(n9063) );
  MUX2X1 U12298 ( .B(n9062), .A(n9059), .S(n10688), .Y(n9073) );
  MUX2X1 U12299 ( .B(\RF[6][17] ), .A(\RF[7][17] ), .S(n10562), .Y(n9067) );
  MUX2X1 U12300 ( .B(\RF[4][17] ), .A(\RF[5][17] ), .S(n10562), .Y(n9066) );
  MUX2X1 U12301 ( .B(\RF[2][17] ), .A(\RF[3][17] ), .S(n10562), .Y(n9070) );
  MUX2X1 U12302 ( .B(\RF[0][17] ), .A(\RF[1][17] ), .S(n10562), .Y(n9069) );
  MUX2X1 U12303 ( .B(n9068), .A(n9065), .S(n10688), .Y(n9072) );
  MUX2X1 U12304 ( .B(n9071), .A(n9056), .S(N22), .Y(n10471) );
  MUX2X1 U12305 ( .B(\RF[30][18] ), .A(\RF[31][18] ), .S(n10562), .Y(n9076) );
  MUX2X1 U12306 ( .B(\RF[28][18] ), .A(\RF[29][18] ), .S(n10562), .Y(n9075) );
  MUX2X1 U12307 ( .B(\RF[26][18] ), .A(\RF[27][18] ), .S(n10562), .Y(n9079) );
  MUX2X1 U12308 ( .B(\RF[24][18] ), .A(\RF[25][18] ), .S(n10562), .Y(n9078) );
  MUX2X1 U12309 ( .B(n9077), .A(n9074), .S(n10688), .Y(n9088) );
  MUX2X1 U12310 ( .B(\RF[22][18] ), .A(\RF[23][18] ), .S(n10563), .Y(n9082) );
  MUX2X1 U12311 ( .B(\RF[20][18] ), .A(\RF[21][18] ), .S(n10563), .Y(n9081) );
  MUX2X1 U12312 ( .B(\RF[18][18] ), .A(\RF[19][18] ), .S(n10563), .Y(n9085) );
  MUX2X1 U12313 ( .B(\RF[16][18] ), .A(\RF[17][18] ), .S(n10563), .Y(n9084) );
  MUX2X1 U12314 ( .B(n9083), .A(n9080), .S(n10688), .Y(n9087) );
  MUX2X1 U12315 ( .B(\RF[14][18] ), .A(\RF[15][18] ), .S(n10563), .Y(n9091) );
  MUX2X1 U12316 ( .B(\RF[12][18] ), .A(\RF[13][18] ), .S(n10563), .Y(n9090) );
  MUX2X1 U12317 ( .B(\RF[10][18] ), .A(\RF[11][18] ), .S(n10563), .Y(n9094) );
  MUX2X1 U12318 ( .B(\RF[8][18] ), .A(\RF[9][18] ), .S(n10563), .Y(n9093) );
  MUX2X1 U12319 ( .B(n9092), .A(n9089), .S(n10688), .Y(n9103) );
  MUX2X1 U12320 ( .B(\RF[6][18] ), .A(\RF[7][18] ), .S(n10563), .Y(n9097) );
  MUX2X1 U12321 ( .B(\RF[4][18] ), .A(\RF[5][18] ), .S(n10563), .Y(n9096) );
  MUX2X1 U12322 ( .B(\RF[2][18] ), .A(\RF[3][18] ), .S(n10563), .Y(n9100) );
  MUX2X1 U12323 ( .B(\RF[0][18] ), .A(\RF[1][18] ), .S(n10563), .Y(n9099) );
  MUX2X1 U12324 ( .B(n9098), .A(n9095), .S(n10688), .Y(n9102) );
  MUX2X1 U12325 ( .B(n9101), .A(n9086), .S(N22), .Y(n10472) );
  MUX2X1 U12326 ( .B(\RF[30][19] ), .A(\RF[31][19] ), .S(n10564), .Y(n9106) );
  MUX2X1 U12327 ( .B(\RF[28][19] ), .A(\RF[29][19] ), .S(n10564), .Y(n9105) );
  MUX2X1 U12328 ( .B(\RF[26][19] ), .A(\RF[27][19] ), .S(n10564), .Y(n9109) );
  MUX2X1 U12329 ( .B(\RF[24][19] ), .A(\RF[25][19] ), .S(n10564), .Y(n9108) );
  MUX2X1 U12330 ( .B(n9107), .A(n9104), .S(n10689), .Y(n9118) );
  MUX2X1 U12331 ( .B(\RF[22][19] ), .A(\RF[23][19] ), .S(n10564), .Y(n9112) );
  MUX2X1 U12332 ( .B(\RF[20][19] ), .A(\RF[21][19] ), .S(n10564), .Y(n9111) );
  MUX2X1 U12333 ( .B(\RF[18][19] ), .A(\RF[19][19] ), .S(n10564), .Y(n9115) );
  MUX2X1 U12334 ( .B(\RF[16][19] ), .A(\RF[17][19] ), .S(n10564), .Y(n9114) );
  MUX2X1 U12335 ( .B(n9113), .A(n9110), .S(n10689), .Y(n9117) );
  MUX2X1 U12336 ( .B(\RF[14][19] ), .A(\RF[15][19] ), .S(n10564), .Y(n9121) );
  MUX2X1 U12337 ( .B(\RF[12][19] ), .A(\RF[13][19] ), .S(n10564), .Y(n9120) );
  MUX2X1 U12338 ( .B(\RF[10][19] ), .A(\RF[11][19] ), .S(n10564), .Y(n9124) );
  MUX2X1 U12339 ( .B(\RF[8][19] ), .A(\RF[9][19] ), .S(n10564), .Y(n9123) );
  MUX2X1 U12340 ( .B(n9122), .A(n9119), .S(n10689), .Y(n9133) );
  MUX2X1 U12341 ( .B(\RF[6][19] ), .A(\RF[7][19] ), .S(n10565), .Y(n9127) );
  MUX2X1 U12342 ( .B(\RF[4][19] ), .A(\RF[5][19] ), .S(n10565), .Y(n9126) );
  MUX2X1 U12343 ( .B(\RF[2][19] ), .A(\RF[3][19] ), .S(n10565), .Y(n9130) );
  MUX2X1 U12344 ( .B(\RF[0][19] ), .A(\RF[1][19] ), .S(n10565), .Y(n9129) );
  MUX2X1 U12345 ( .B(n9128), .A(n9125), .S(n10689), .Y(n9132) );
  MUX2X1 U12346 ( .B(n9131), .A(n9116), .S(N22), .Y(n10473) );
  MUX2X1 U12347 ( .B(\RF[30][20] ), .A(\RF[31][20] ), .S(n10565), .Y(n9136) );
  MUX2X1 U12348 ( .B(\RF[28][20] ), .A(\RF[29][20] ), .S(n10565), .Y(n9135) );
  MUX2X1 U12349 ( .B(\RF[26][20] ), .A(\RF[27][20] ), .S(n10565), .Y(n9139) );
  MUX2X1 U12350 ( .B(\RF[24][20] ), .A(\RF[25][20] ), .S(n10565), .Y(n9138) );
  MUX2X1 U12351 ( .B(n9137), .A(n9134), .S(n10689), .Y(n9148) );
  MUX2X1 U12352 ( .B(\RF[22][20] ), .A(\RF[23][20] ), .S(n10565), .Y(n9142) );
  MUX2X1 U12353 ( .B(\RF[20][20] ), .A(\RF[21][20] ), .S(n10565), .Y(n9141) );
  MUX2X1 U12354 ( .B(\RF[18][20] ), .A(\RF[19][20] ), .S(n10565), .Y(n9145) );
  MUX2X1 U12355 ( .B(\RF[16][20] ), .A(\RF[17][20] ), .S(n10565), .Y(n9144) );
  MUX2X1 U12356 ( .B(n9143), .A(n9140), .S(n10689), .Y(n9147) );
  MUX2X1 U12357 ( .B(\RF[14][20] ), .A(\RF[15][20] ), .S(n10566), .Y(n9151) );
  MUX2X1 U12358 ( .B(\RF[12][20] ), .A(\RF[13][20] ), .S(n10566), .Y(n9150) );
  MUX2X1 U12359 ( .B(\RF[10][20] ), .A(\RF[11][20] ), .S(n10566), .Y(n9154) );
  MUX2X1 U12360 ( .B(\RF[8][20] ), .A(\RF[9][20] ), .S(n10566), .Y(n9153) );
  MUX2X1 U12361 ( .B(n9152), .A(n9149), .S(n10689), .Y(n9163) );
  MUX2X1 U12362 ( .B(\RF[6][20] ), .A(\RF[7][20] ), .S(n10566), .Y(n9157) );
  MUX2X1 U12363 ( .B(\RF[4][20] ), .A(\RF[5][20] ), .S(n10566), .Y(n9156) );
  MUX2X1 U12364 ( .B(\RF[2][20] ), .A(\RF[3][20] ), .S(n10566), .Y(n9160) );
  MUX2X1 U12365 ( .B(\RF[0][20] ), .A(\RF[1][20] ), .S(n10566), .Y(n9159) );
  MUX2X1 U12366 ( .B(n9158), .A(n9155), .S(n10689), .Y(n9162) );
  MUX2X1 U12367 ( .B(n9161), .A(n9146), .S(N22), .Y(n10474) );
  MUX2X1 U12368 ( .B(\RF[30][21] ), .A(\RF[31][21] ), .S(n10566), .Y(n9166) );
  MUX2X1 U12369 ( .B(\RF[28][21] ), .A(\RF[29][21] ), .S(n10566), .Y(n9165) );
  MUX2X1 U12370 ( .B(\RF[26][21] ), .A(\RF[27][21] ), .S(n10566), .Y(n9169) );
  MUX2X1 U12371 ( .B(\RF[24][21] ), .A(\RF[25][21] ), .S(n10566), .Y(n9168) );
  MUX2X1 U12372 ( .B(n9167), .A(n9164), .S(n10689), .Y(n9178) );
  MUX2X1 U12373 ( .B(\RF[22][21] ), .A(\RF[23][21] ), .S(n10567), .Y(n9172) );
  MUX2X1 U12374 ( .B(\RF[20][21] ), .A(\RF[21][21] ), .S(n10567), .Y(n9171) );
  MUX2X1 U12375 ( .B(\RF[18][21] ), .A(\RF[19][21] ), .S(n10567), .Y(n9175) );
  MUX2X1 U12376 ( .B(\RF[16][21] ), .A(\RF[17][21] ), .S(n10567), .Y(n9174) );
  MUX2X1 U12377 ( .B(n9173), .A(n9170), .S(n10689), .Y(n9177) );
  MUX2X1 U12378 ( .B(\RF[14][21] ), .A(\RF[15][21] ), .S(n10567), .Y(n9181) );
  MUX2X1 U12379 ( .B(\RF[12][21] ), .A(\RF[13][21] ), .S(n10567), .Y(n9180) );
  MUX2X1 U12380 ( .B(\RF[10][21] ), .A(\RF[11][21] ), .S(n10567), .Y(n9184) );
  MUX2X1 U12381 ( .B(\RF[8][21] ), .A(\RF[9][21] ), .S(n10567), .Y(n9183) );
  MUX2X1 U12382 ( .B(n9182), .A(n9179), .S(n10689), .Y(n9193) );
  MUX2X1 U12383 ( .B(\RF[6][21] ), .A(\RF[7][21] ), .S(n10567), .Y(n9187) );
  MUX2X1 U12384 ( .B(\RF[4][21] ), .A(\RF[5][21] ), .S(n10567), .Y(n9186) );
  MUX2X1 U12385 ( .B(\RF[2][21] ), .A(\RF[3][21] ), .S(n10567), .Y(n9190) );
  MUX2X1 U12386 ( .B(\RF[0][21] ), .A(\RF[1][21] ), .S(n10567), .Y(n9189) );
  MUX2X1 U12387 ( .B(n9188), .A(n9185), .S(n10689), .Y(n9192) );
  MUX2X1 U12388 ( .B(n9191), .A(n9176), .S(N22), .Y(n10475) );
  MUX2X1 U12389 ( .B(\RF[30][22] ), .A(\RF[31][22] ), .S(n10568), .Y(n9196) );
  MUX2X1 U12390 ( .B(\RF[28][22] ), .A(\RF[29][22] ), .S(n10568), .Y(n9195) );
  MUX2X1 U12391 ( .B(\RF[26][22] ), .A(\RF[27][22] ), .S(n10568), .Y(n9199) );
  MUX2X1 U12392 ( .B(\RF[24][22] ), .A(\RF[25][22] ), .S(n10568), .Y(n9198) );
  MUX2X1 U12393 ( .B(n9197), .A(n9194), .S(n10690), .Y(n9208) );
  MUX2X1 U12394 ( .B(\RF[22][22] ), .A(\RF[23][22] ), .S(n10568), .Y(n9202) );
  MUX2X1 U12395 ( .B(\RF[20][22] ), .A(\RF[21][22] ), .S(n10568), .Y(n9201) );
  MUX2X1 U12396 ( .B(\RF[18][22] ), .A(\RF[19][22] ), .S(n10568), .Y(n9205) );
  MUX2X1 U12397 ( .B(\RF[16][22] ), .A(\RF[17][22] ), .S(n10568), .Y(n9204) );
  MUX2X1 U12398 ( .B(n9203), .A(n9200), .S(n10690), .Y(n9207) );
  MUX2X1 U12399 ( .B(\RF[14][22] ), .A(\RF[15][22] ), .S(n10568), .Y(n9211) );
  MUX2X1 U12400 ( .B(\RF[12][22] ), .A(\RF[13][22] ), .S(n10568), .Y(n9210) );
  MUX2X1 U12401 ( .B(\RF[10][22] ), .A(\RF[11][22] ), .S(n10568), .Y(n9214) );
  MUX2X1 U12402 ( .B(\RF[8][22] ), .A(\RF[9][22] ), .S(n10568), .Y(n9213) );
  MUX2X1 U12403 ( .B(n9212), .A(n9209), .S(n10690), .Y(n9223) );
  MUX2X1 U12404 ( .B(\RF[6][22] ), .A(\RF[7][22] ), .S(n10569), .Y(n9217) );
  MUX2X1 U12405 ( .B(\RF[4][22] ), .A(\RF[5][22] ), .S(n10569), .Y(n9216) );
  MUX2X1 U12406 ( .B(\RF[2][22] ), .A(\RF[3][22] ), .S(n10569), .Y(n9220) );
  MUX2X1 U12407 ( .B(\RF[0][22] ), .A(\RF[1][22] ), .S(n10569), .Y(n9219) );
  MUX2X1 U12408 ( .B(n9218), .A(n9215), .S(n10690), .Y(n9222) );
  MUX2X1 U12409 ( .B(n9221), .A(n9206), .S(N22), .Y(n10476) );
  MUX2X1 U12410 ( .B(\RF[30][23] ), .A(\RF[31][23] ), .S(n10569), .Y(n9226) );
  MUX2X1 U12411 ( .B(\RF[28][23] ), .A(\RF[29][23] ), .S(n10569), .Y(n9225) );
  MUX2X1 U12412 ( .B(\RF[26][23] ), .A(\RF[27][23] ), .S(n10569), .Y(n9229) );
  MUX2X1 U12413 ( .B(\RF[24][23] ), .A(\RF[25][23] ), .S(n10569), .Y(n9228) );
  MUX2X1 U12414 ( .B(n9227), .A(n9224), .S(n10690), .Y(n9238) );
  MUX2X1 U12415 ( .B(\RF[22][23] ), .A(\RF[23][23] ), .S(n10569), .Y(n9232) );
  MUX2X1 U12416 ( .B(\RF[20][23] ), .A(\RF[21][23] ), .S(n10569), .Y(n9231) );
  MUX2X1 U12417 ( .B(\RF[18][23] ), .A(\RF[19][23] ), .S(n10569), .Y(n9235) );
  MUX2X1 U12418 ( .B(\RF[16][23] ), .A(\RF[17][23] ), .S(n10569), .Y(n9234) );
  MUX2X1 U12419 ( .B(n9233), .A(n9230), .S(n10690), .Y(n9237) );
  MUX2X1 U12420 ( .B(\RF[14][23] ), .A(\RF[15][23] ), .S(n10570), .Y(n9241) );
  MUX2X1 U12421 ( .B(\RF[12][23] ), .A(\RF[13][23] ), .S(n10570), .Y(n9240) );
  MUX2X1 U12422 ( .B(\RF[10][23] ), .A(\RF[11][23] ), .S(n10570), .Y(n9244) );
  MUX2X1 U12423 ( .B(\RF[8][23] ), .A(\RF[9][23] ), .S(n10570), .Y(n9243) );
  MUX2X1 U12424 ( .B(n9242), .A(n9239), .S(n10690), .Y(n9253) );
  MUX2X1 U12425 ( .B(\RF[6][23] ), .A(\RF[7][23] ), .S(n10570), .Y(n9247) );
  MUX2X1 U12426 ( .B(\RF[4][23] ), .A(\RF[5][23] ), .S(n10570), .Y(n9246) );
  MUX2X1 U12427 ( .B(\RF[2][23] ), .A(\RF[3][23] ), .S(n10570), .Y(n9250) );
  MUX2X1 U12428 ( .B(\RF[0][23] ), .A(\RF[1][23] ), .S(n10570), .Y(n9249) );
  MUX2X1 U12429 ( .B(n9248), .A(n9245), .S(n10690), .Y(n9252) );
  MUX2X1 U12430 ( .B(n9251), .A(n9236), .S(N22), .Y(n10477) );
  MUX2X1 U12431 ( .B(\RF[30][24] ), .A(\RF[31][24] ), .S(n10570), .Y(n9256) );
  MUX2X1 U12432 ( .B(\RF[28][24] ), .A(\RF[29][24] ), .S(n10570), .Y(n9255) );
  MUX2X1 U12433 ( .B(\RF[26][24] ), .A(\RF[27][24] ), .S(n10570), .Y(n9259) );
  MUX2X1 U12434 ( .B(\RF[24][24] ), .A(\RF[25][24] ), .S(n10570), .Y(n9258) );
  MUX2X1 U12435 ( .B(n9257), .A(n9254), .S(n10690), .Y(n9268) );
  MUX2X1 U12436 ( .B(\RF[22][24] ), .A(\RF[23][24] ), .S(n10571), .Y(n9262) );
  MUX2X1 U12437 ( .B(\RF[20][24] ), .A(\RF[21][24] ), .S(n10571), .Y(n9261) );
  MUX2X1 U12438 ( .B(\RF[18][24] ), .A(\RF[19][24] ), .S(n10571), .Y(n9265) );
  MUX2X1 U12439 ( .B(\RF[16][24] ), .A(\RF[17][24] ), .S(n10571), .Y(n9264) );
  MUX2X1 U12440 ( .B(n9263), .A(n9260), .S(n10690), .Y(n9267) );
  MUX2X1 U12441 ( .B(\RF[14][24] ), .A(\RF[15][24] ), .S(n10571), .Y(n9271) );
  MUX2X1 U12442 ( .B(\RF[12][24] ), .A(\RF[13][24] ), .S(n10571), .Y(n9270) );
  MUX2X1 U12443 ( .B(\RF[10][24] ), .A(\RF[11][24] ), .S(n10571), .Y(n9274) );
  MUX2X1 U12444 ( .B(\RF[8][24] ), .A(\RF[9][24] ), .S(n10571), .Y(n9273) );
  MUX2X1 U12445 ( .B(n9272), .A(n9269), .S(n10690), .Y(n9283) );
  MUX2X1 U12446 ( .B(\RF[6][24] ), .A(\RF[7][24] ), .S(n10571), .Y(n9277) );
  MUX2X1 U12447 ( .B(\RF[4][24] ), .A(\RF[5][24] ), .S(n10571), .Y(n9276) );
  MUX2X1 U12448 ( .B(\RF[2][24] ), .A(\RF[3][24] ), .S(n10571), .Y(n9280) );
  MUX2X1 U12449 ( .B(\RF[0][24] ), .A(\RF[1][24] ), .S(n10571), .Y(n9279) );
  MUX2X1 U12450 ( .B(n9278), .A(n9275), .S(n10690), .Y(n9282) );
  MUX2X1 U12451 ( .B(n9281), .A(n9266), .S(N22), .Y(n10478) );
  MUX2X1 U12452 ( .B(\RF[30][25] ), .A(\RF[31][25] ), .S(n10572), .Y(n9286) );
  MUX2X1 U12453 ( .B(\RF[28][25] ), .A(\RF[29][25] ), .S(n10572), .Y(n9285) );
  MUX2X1 U12454 ( .B(\RF[26][25] ), .A(\RF[27][25] ), .S(n10572), .Y(n9289) );
  MUX2X1 U12455 ( .B(\RF[24][25] ), .A(\RF[25][25] ), .S(n10572), .Y(n9288) );
  MUX2X1 U12456 ( .B(n9287), .A(n9284), .S(n10691), .Y(n9298) );
  MUX2X1 U12457 ( .B(\RF[22][25] ), .A(\RF[23][25] ), .S(n10572), .Y(n9292) );
  MUX2X1 U12458 ( .B(\RF[20][25] ), .A(\RF[21][25] ), .S(n10572), .Y(n9291) );
  MUX2X1 U12459 ( .B(\RF[18][25] ), .A(\RF[19][25] ), .S(n10572), .Y(n9295) );
  MUX2X1 U12460 ( .B(\RF[16][25] ), .A(\RF[17][25] ), .S(n10572), .Y(n9294) );
  MUX2X1 U12461 ( .B(n9293), .A(n9290), .S(n10691), .Y(n9297) );
  MUX2X1 U12462 ( .B(\RF[14][25] ), .A(\RF[15][25] ), .S(n10572), .Y(n9301) );
  MUX2X1 U12463 ( .B(\RF[12][25] ), .A(\RF[13][25] ), .S(n10572), .Y(n9300) );
  MUX2X1 U12464 ( .B(\RF[10][25] ), .A(\RF[11][25] ), .S(n10572), .Y(n9304) );
  MUX2X1 U12465 ( .B(\RF[8][25] ), .A(\RF[9][25] ), .S(n10572), .Y(n9303) );
  MUX2X1 U12466 ( .B(n9302), .A(n9299), .S(n10691), .Y(n9313) );
  MUX2X1 U12467 ( .B(\RF[6][25] ), .A(\RF[7][25] ), .S(n10573), .Y(n9307) );
  MUX2X1 U12468 ( .B(\RF[4][25] ), .A(\RF[5][25] ), .S(n10573), .Y(n9306) );
  MUX2X1 U12469 ( .B(\RF[2][25] ), .A(\RF[3][25] ), .S(n10573), .Y(n9310) );
  MUX2X1 U12470 ( .B(\RF[0][25] ), .A(\RF[1][25] ), .S(n10573), .Y(n9309) );
  MUX2X1 U12471 ( .B(n9308), .A(n9305), .S(n10691), .Y(n9312) );
  MUX2X1 U12472 ( .B(n9311), .A(n9296), .S(N22), .Y(n10479) );
  MUX2X1 U12473 ( .B(\RF[30][26] ), .A(\RF[31][26] ), .S(n10573), .Y(n9316) );
  MUX2X1 U12474 ( .B(\RF[28][26] ), .A(\RF[29][26] ), .S(n10573), .Y(n9315) );
  MUX2X1 U12475 ( .B(\RF[26][26] ), .A(\RF[27][26] ), .S(n10573), .Y(n9319) );
  MUX2X1 U12476 ( .B(\RF[24][26] ), .A(\RF[25][26] ), .S(n10573), .Y(n9318) );
  MUX2X1 U12477 ( .B(n9317), .A(n9314), .S(n10691), .Y(n9328) );
  MUX2X1 U12478 ( .B(\RF[22][26] ), .A(\RF[23][26] ), .S(n10573), .Y(n9322) );
  MUX2X1 U12479 ( .B(\RF[20][26] ), .A(\RF[21][26] ), .S(n10573), .Y(n9321) );
  MUX2X1 U12480 ( .B(\RF[18][26] ), .A(\RF[19][26] ), .S(n10573), .Y(n9325) );
  MUX2X1 U12481 ( .B(\RF[16][26] ), .A(\RF[17][26] ), .S(n10573), .Y(n9324) );
  MUX2X1 U12482 ( .B(n9323), .A(n9320), .S(n10691), .Y(n9327) );
  MUX2X1 U12483 ( .B(\RF[14][26] ), .A(\RF[15][26] ), .S(n10574), .Y(n9331) );
  MUX2X1 U12484 ( .B(\RF[12][26] ), .A(\RF[13][26] ), .S(n10574), .Y(n9330) );
  MUX2X1 U12485 ( .B(\RF[10][26] ), .A(\RF[11][26] ), .S(n10574), .Y(n9334) );
  MUX2X1 U12486 ( .B(\RF[8][26] ), .A(\RF[9][26] ), .S(n10574), .Y(n9333) );
  MUX2X1 U12487 ( .B(n9332), .A(n9329), .S(n10691), .Y(n9343) );
  MUX2X1 U12488 ( .B(\RF[6][26] ), .A(\RF[7][26] ), .S(n10574), .Y(n9337) );
  MUX2X1 U12489 ( .B(\RF[4][26] ), .A(\RF[5][26] ), .S(n10574), .Y(n9336) );
  MUX2X1 U12490 ( .B(\RF[2][26] ), .A(\RF[3][26] ), .S(n10574), .Y(n9340) );
  MUX2X1 U12491 ( .B(\RF[0][26] ), .A(\RF[1][26] ), .S(n10574), .Y(n9339) );
  MUX2X1 U12492 ( .B(n9338), .A(n9335), .S(n10691), .Y(n9342) );
  MUX2X1 U12493 ( .B(n9341), .A(n9326), .S(N22), .Y(n10480) );
  MUX2X1 U12494 ( .B(\RF[30][27] ), .A(\RF[31][27] ), .S(n10574), .Y(n9346) );
  MUX2X1 U12495 ( .B(\RF[28][27] ), .A(\RF[29][27] ), .S(n10574), .Y(n9345) );
  MUX2X1 U12496 ( .B(\RF[26][27] ), .A(\RF[27][27] ), .S(n10574), .Y(n9349) );
  MUX2X1 U12497 ( .B(\RF[24][27] ), .A(\RF[25][27] ), .S(n10574), .Y(n9348) );
  MUX2X1 U12498 ( .B(n9347), .A(n9344), .S(n10691), .Y(n9358) );
  MUX2X1 U12499 ( .B(\RF[22][27] ), .A(\RF[23][27] ), .S(n10575), .Y(n9352) );
  MUX2X1 U12500 ( .B(\RF[20][27] ), .A(\RF[21][27] ), .S(n10575), .Y(n9351) );
  MUX2X1 U12501 ( .B(\RF[18][27] ), .A(\RF[19][27] ), .S(n10575), .Y(n9355) );
  MUX2X1 U12502 ( .B(\RF[16][27] ), .A(\RF[17][27] ), .S(n10575), .Y(n9354) );
  MUX2X1 U12503 ( .B(n9353), .A(n9350), .S(n10691), .Y(n9357) );
  MUX2X1 U12504 ( .B(\RF[14][27] ), .A(\RF[15][27] ), .S(n10575), .Y(n9361) );
  MUX2X1 U12505 ( .B(\RF[12][27] ), .A(\RF[13][27] ), .S(n10575), .Y(n9360) );
  MUX2X1 U12506 ( .B(\RF[10][27] ), .A(\RF[11][27] ), .S(n10575), .Y(n9364) );
  MUX2X1 U12507 ( .B(\RF[8][27] ), .A(\RF[9][27] ), .S(n10575), .Y(n9363) );
  MUX2X1 U12508 ( .B(n9362), .A(n9359), .S(n10691), .Y(n9373) );
  MUX2X1 U12509 ( .B(\RF[6][27] ), .A(\RF[7][27] ), .S(n10575), .Y(n9367) );
  MUX2X1 U12510 ( .B(\RF[4][27] ), .A(\RF[5][27] ), .S(n10575), .Y(n9366) );
  MUX2X1 U12511 ( .B(\RF[2][27] ), .A(\RF[3][27] ), .S(n10575), .Y(n9370) );
  MUX2X1 U12512 ( .B(\RF[0][27] ), .A(\RF[1][27] ), .S(n10575), .Y(n9369) );
  MUX2X1 U12513 ( .B(n9368), .A(n9365), .S(n10691), .Y(n9372) );
  MUX2X1 U12514 ( .B(n9371), .A(n9356), .S(N22), .Y(n10481) );
  MUX2X1 U12515 ( .B(\RF[30][28] ), .A(\RF[31][28] ), .S(n10576), .Y(n9376) );
  MUX2X1 U12516 ( .B(\RF[28][28] ), .A(\RF[29][28] ), .S(n10576), .Y(n9375) );
  MUX2X1 U12517 ( .B(\RF[26][28] ), .A(\RF[27][28] ), .S(n10576), .Y(n9379) );
  MUX2X1 U12518 ( .B(\RF[24][28] ), .A(\RF[25][28] ), .S(n10576), .Y(n9378) );
  MUX2X1 U12519 ( .B(n9377), .A(n9374), .S(n10692), .Y(n9388) );
  MUX2X1 U12520 ( .B(\RF[22][28] ), .A(\RF[23][28] ), .S(n10576), .Y(n9382) );
  MUX2X1 U12521 ( .B(\RF[20][28] ), .A(\RF[21][28] ), .S(n10576), .Y(n9381) );
  MUX2X1 U12522 ( .B(\RF[18][28] ), .A(\RF[19][28] ), .S(n10576), .Y(n9385) );
  MUX2X1 U12523 ( .B(\RF[16][28] ), .A(\RF[17][28] ), .S(n10576), .Y(n9384) );
  MUX2X1 U12524 ( .B(n9383), .A(n9380), .S(n10692), .Y(n9387) );
  MUX2X1 U12525 ( .B(\RF[14][28] ), .A(\RF[15][28] ), .S(n10576), .Y(n9391) );
  MUX2X1 U12526 ( .B(\RF[12][28] ), .A(\RF[13][28] ), .S(n10576), .Y(n9390) );
  MUX2X1 U12527 ( .B(\RF[10][28] ), .A(\RF[11][28] ), .S(n10576), .Y(n9394) );
  MUX2X1 U12528 ( .B(\RF[8][28] ), .A(\RF[9][28] ), .S(n10576), .Y(n9393) );
  MUX2X1 U12529 ( .B(n9392), .A(n9389), .S(n10692), .Y(n9403) );
  MUX2X1 U12530 ( .B(\RF[6][28] ), .A(\RF[7][28] ), .S(n10577), .Y(n9397) );
  MUX2X1 U12531 ( .B(\RF[4][28] ), .A(\RF[5][28] ), .S(n10577), .Y(n9396) );
  MUX2X1 U12532 ( .B(\RF[2][28] ), .A(\RF[3][28] ), .S(n10577), .Y(n9400) );
  MUX2X1 U12533 ( .B(\RF[0][28] ), .A(\RF[1][28] ), .S(n10577), .Y(n9399) );
  MUX2X1 U12534 ( .B(n9398), .A(n9395), .S(n10692), .Y(n9402) );
  MUX2X1 U12535 ( .B(n9401), .A(n9386), .S(N22), .Y(n10482) );
  MUX2X1 U12536 ( .B(\RF[30][29] ), .A(\RF[31][29] ), .S(n10577), .Y(n9406) );
  MUX2X1 U12537 ( .B(\RF[28][29] ), .A(\RF[29][29] ), .S(n10577), .Y(n9405) );
  MUX2X1 U12538 ( .B(\RF[26][29] ), .A(\RF[27][29] ), .S(n10577), .Y(n9409) );
  MUX2X1 U12539 ( .B(\RF[24][29] ), .A(\RF[25][29] ), .S(n10577), .Y(n9408) );
  MUX2X1 U12540 ( .B(n9407), .A(n9404), .S(n10692), .Y(n9418) );
  MUX2X1 U12541 ( .B(\RF[22][29] ), .A(\RF[23][29] ), .S(n10577), .Y(n9412) );
  MUX2X1 U12542 ( .B(\RF[20][29] ), .A(\RF[21][29] ), .S(n10577), .Y(n9411) );
  MUX2X1 U12543 ( .B(\RF[18][29] ), .A(\RF[19][29] ), .S(n10577), .Y(n9415) );
  MUX2X1 U12544 ( .B(\RF[16][29] ), .A(\RF[17][29] ), .S(n10577), .Y(n9414) );
  MUX2X1 U12545 ( .B(n9413), .A(n9410), .S(n10692), .Y(n9417) );
  MUX2X1 U12546 ( .B(\RF[14][29] ), .A(\RF[15][29] ), .S(n10578), .Y(n9421) );
  MUX2X1 U12547 ( .B(\RF[12][29] ), .A(\RF[13][29] ), .S(n10578), .Y(n9420) );
  MUX2X1 U12548 ( .B(\RF[10][29] ), .A(\RF[11][29] ), .S(n10578), .Y(n9424) );
  MUX2X1 U12549 ( .B(\RF[8][29] ), .A(\RF[9][29] ), .S(n10578), .Y(n9423) );
  MUX2X1 U12550 ( .B(n9422), .A(n9419), .S(n10692), .Y(n9433) );
  MUX2X1 U12551 ( .B(\RF[6][29] ), .A(\RF[7][29] ), .S(n10578), .Y(n9427) );
  MUX2X1 U12552 ( .B(\RF[4][29] ), .A(\RF[5][29] ), .S(n10578), .Y(n9426) );
  MUX2X1 U12553 ( .B(\RF[2][29] ), .A(\RF[3][29] ), .S(n10578), .Y(n9430) );
  MUX2X1 U12554 ( .B(\RF[0][29] ), .A(\RF[1][29] ), .S(n10578), .Y(n9429) );
  MUX2X1 U12555 ( .B(n9428), .A(n9425), .S(n10692), .Y(n9432) );
  MUX2X1 U12556 ( .B(n9431), .A(n9416), .S(N22), .Y(n10483) );
  MUX2X1 U12557 ( .B(\RF[30][30] ), .A(\RF[31][30] ), .S(n10578), .Y(n9436) );
  MUX2X1 U12558 ( .B(\RF[28][30] ), .A(\RF[29][30] ), .S(n10578), .Y(n9435) );
  MUX2X1 U12559 ( .B(\RF[26][30] ), .A(\RF[27][30] ), .S(n10578), .Y(n9439) );
  MUX2X1 U12560 ( .B(\RF[24][30] ), .A(\RF[25][30] ), .S(n10578), .Y(n9438) );
  MUX2X1 U12561 ( .B(n9437), .A(n9434), .S(n10692), .Y(n9448) );
  MUX2X1 U12562 ( .B(\RF[22][30] ), .A(\RF[23][30] ), .S(n10579), .Y(n9442) );
  MUX2X1 U12563 ( .B(\RF[20][30] ), .A(\RF[21][30] ), .S(n10579), .Y(n9441) );
  MUX2X1 U12564 ( .B(\RF[18][30] ), .A(\RF[19][30] ), .S(n10579), .Y(n9445) );
  MUX2X1 U12565 ( .B(\RF[16][30] ), .A(\RF[17][30] ), .S(n10579), .Y(n9444) );
  MUX2X1 U12566 ( .B(n9443), .A(n9440), .S(n10692), .Y(n9447) );
  MUX2X1 U12567 ( .B(\RF[14][30] ), .A(\RF[15][30] ), .S(n10579), .Y(n9451) );
  MUX2X1 U12568 ( .B(\RF[12][30] ), .A(\RF[13][30] ), .S(n10579), .Y(n9450) );
  MUX2X1 U12569 ( .B(\RF[10][30] ), .A(\RF[11][30] ), .S(n10579), .Y(n9454) );
  MUX2X1 U12570 ( .B(\RF[8][30] ), .A(\RF[9][30] ), .S(n10579), .Y(n9453) );
  MUX2X1 U12571 ( .B(n9452), .A(n9449), .S(n10692), .Y(n9463) );
  MUX2X1 U12572 ( .B(\RF[6][30] ), .A(\RF[7][30] ), .S(n10579), .Y(n9457) );
  MUX2X1 U12573 ( .B(\RF[4][30] ), .A(\RF[5][30] ), .S(n10579), .Y(n9456) );
  MUX2X1 U12574 ( .B(\RF[2][30] ), .A(\RF[3][30] ), .S(n10579), .Y(n9460) );
  MUX2X1 U12575 ( .B(\RF[0][30] ), .A(\RF[1][30] ), .S(n10579), .Y(n9459) );
  MUX2X1 U12576 ( .B(n9458), .A(n9455), .S(n10692), .Y(n9462) );
  MUX2X1 U12577 ( .B(n9461), .A(n9446), .S(N22), .Y(n10484) );
  MUX2X1 U12578 ( .B(\RF[30][31] ), .A(\RF[31][31] ), .S(n10580), .Y(n9466) );
  MUX2X1 U12579 ( .B(\RF[28][31] ), .A(\RF[29][31] ), .S(n10580), .Y(n9465) );
  MUX2X1 U12580 ( .B(\RF[26][31] ), .A(\RF[27][31] ), .S(n10580), .Y(n9469) );
  MUX2X1 U12581 ( .B(\RF[24][31] ), .A(\RF[25][31] ), .S(n10580), .Y(n9468) );
  MUX2X1 U12582 ( .B(n9467), .A(n9464), .S(n10693), .Y(n9478) );
  MUX2X1 U12583 ( .B(\RF[22][31] ), .A(\RF[23][31] ), .S(n10580), .Y(n9472) );
  MUX2X1 U12584 ( .B(\RF[20][31] ), .A(\RF[21][31] ), .S(n10580), .Y(n9471) );
  MUX2X1 U12585 ( .B(\RF[18][31] ), .A(\RF[19][31] ), .S(n10580), .Y(n9475) );
  MUX2X1 U12586 ( .B(\RF[16][31] ), .A(\RF[17][31] ), .S(n10580), .Y(n9474) );
  MUX2X1 U12587 ( .B(n9473), .A(n9470), .S(n10693), .Y(n9477) );
  MUX2X1 U12588 ( .B(\RF[14][31] ), .A(\RF[15][31] ), .S(n10580), .Y(n9481) );
  MUX2X1 U12589 ( .B(\RF[12][31] ), .A(\RF[13][31] ), .S(n10580), .Y(n9480) );
  MUX2X1 U12590 ( .B(\RF[10][31] ), .A(\RF[11][31] ), .S(n10580), .Y(n9484) );
  MUX2X1 U12591 ( .B(\RF[8][31] ), .A(\RF[9][31] ), .S(n10580), .Y(n9483) );
  MUX2X1 U12592 ( .B(n9482), .A(n9479), .S(n10693), .Y(n9493) );
  MUX2X1 U12593 ( .B(\RF[6][31] ), .A(\RF[7][31] ), .S(n10581), .Y(n9487) );
  MUX2X1 U12594 ( .B(\RF[4][31] ), .A(\RF[5][31] ), .S(n10581), .Y(n9486) );
  MUX2X1 U12595 ( .B(\RF[2][31] ), .A(\RF[3][31] ), .S(n10581), .Y(n9490) );
  MUX2X1 U12596 ( .B(\RF[0][31] ), .A(\RF[1][31] ), .S(n10581), .Y(n9489) );
  MUX2X1 U12597 ( .B(n9488), .A(n9485), .S(n10693), .Y(n9492) );
  MUX2X1 U12598 ( .B(n9491), .A(n9476), .S(N22), .Y(n10485) );
  MUX2X1 U12599 ( .B(\RF[30][32] ), .A(\RF[31][32] ), .S(n10581), .Y(n9496) );
  MUX2X1 U12600 ( .B(\RF[28][32] ), .A(\RF[29][32] ), .S(n10581), .Y(n9495) );
  MUX2X1 U12601 ( .B(\RF[26][32] ), .A(\RF[27][32] ), .S(n10581), .Y(n9499) );
  MUX2X1 U12602 ( .B(\RF[24][32] ), .A(\RF[25][32] ), .S(n10581), .Y(n9498) );
  MUX2X1 U12603 ( .B(n9497), .A(n9494), .S(n10693), .Y(n9508) );
  MUX2X1 U12604 ( .B(\RF[22][32] ), .A(\RF[23][32] ), .S(n10581), .Y(n9502) );
  MUX2X1 U12605 ( .B(\RF[20][32] ), .A(\RF[21][32] ), .S(n10581), .Y(n9501) );
  MUX2X1 U12606 ( .B(\RF[18][32] ), .A(\RF[19][32] ), .S(n10581), .Y(n9505) );
  MUX2X1 U12607 ( .B(\RF[16][32] ), .A(\RF[17][32] ), .S(n10581), .Y(n9504) );
  MUX2X1 U12608 ( .B(n9503), .A(n9500), .S(n10693), .Y(n9507) );
  MUX2X1 U12609 ( .B(\RF[14][32] ), .A(\RF[15][32] ), .S(n10582), .Y(n9511) );
  MUX2X1 U12610 ( .B(\RF[12][32] ), .A(\RF[13][32] ), .S(n10582), .Y(n9510) );
  MUX2X1 U12611 ( .B(\RF[10][32] ), .A(\RF[11][32] ), .S(n10582), .Y(n9514) );
  MUX2X1 U12612 ( .B(\RF[8][32] ), .A(\RF[9][32] ), .S(n10582), .Y(n9513) );
  MUX2X1 U12613 ( .B(n9512), .A(n9509), .S(n10693), .Y(n9523) );
  MUX2X1 U12614 ( .B(\RF[6][32] ), .A(\RF[7][32] ), .S(n10582), .Y(n9517) );
  MUX2X1 U12615 ( .B(\RF[4][32] ), .A(\RF[5][32] ), .S(n10582), .Y(n9516) );
  MUX2X1 U12616 ( .B(\RF[2][32] ), .A(\RF[3][32] ), .S(n10582), .Y(n9520) );
  MUX2X1 U12617 ( .B(\RF[0][32] ), .A(\RF[1][32] ), .S(n10582), .Y(n9519) );
  MUX2X1 U12618 ( .B(n9518), .A(n9515), .S(n10693), .Y(n9522) );
  MUX2X1 U12619 ( .B(n9521), .A(n9506), .S(N22), .Y(n10486) );
  MUX2X1 U12620 ( .B(\RF[30][33] ), .A(\RF[31][33] ), .S(n10582), .Y(n9526) );
  MUX2X1 U12621 ( .B(\RF[28][33] ), .A(\RF[29][33] ), .S(n10582), .Y(n9525) );
  MUX2X1 U12622 ( .B(\RF[26][33] ), .A(\RF[27][33] ), .S(n10582), .Y(n9529) );
  MUX2X1 U12623 ( .B(\RF[24][33] ), .A(\RF[25][33] ), .S(n10582), .Y(n9528) );
  MUX2X1 U12624 ( .B(n9527), .A(n9524), .S(n10693), .Y(n9538) );
  MUX2X1 U12625 ( .B(\RF[22][33] ), .A(\RF[23][33] ), .S(n10583), .Y(n9532) );
  MUX2X1 U12626 ( .B(\RF[20][33] ), .A(\RF[21][33] ), .S(n10583), .Y(n9531) );
  MUX2X1 U12627 ( .B(\RF[18][33] ), .A(\RF[19][33] ), .S(n10583), .Y(n9535) );
  MUX2X1 U12628 ( .B(\RF[16][33] ), .A(\RF[17][33] ), .S(n10583), .Y(n9534) );
  MUX2X1 U12629 ( .B(n9533), .A(n9530), .S(n10693), .Y(n9537) );
  MUX2X1 U12630 ( .B(\RF[14][33] ), .A(\RF[15][33] ), .S(n10583), .Y(n9541) );
  MUX2X1 U12631 ( .B(\RF[12][33] ), .A(\RF[13][33] ), .S(n10583), .Y(n9540) );
  MUX2X1 U12632 ( .B(\RF[10][33] ), .A(\RF[11][33] ), .S(n10583), .Y(n9544) );
  MUX2X1 U12633 ( .B(\RF[8][33] ), .A(\RF[9][33] ), .S(n10583), .Y(n9543) );
  MUX2X1 U12634 ( .B(n9542), .A(n9539), .S(n10693), .Y(n9553) );
  MUX2X1 U12635 ( .B(\RF[6][33] ), .A(\RF[7][33] ), .S(n10583), .Y(n9547) );
  MUX2X1 U12636 ( .B(\RF[4][33] ), .A(\RF[5][33] ), .S(n10583), .Y(n9546) );
  MUX2X1 U12637 ( .B(\RF[2][33] ), .A(\RF[3][33] ), .S(n10583), .Y(n9550) );
  MUX2X1 U12638 ( .B(\RF[0][33] ), .A(\RF[1][33] ), .S(n10583), .Y(n9549) );
  MUX2X1 U12639 ( .B(n9548), .A(n9545), .S(n10693), .Y(n9552) );
  MUX2X1 U12640 ( .B(n9551), .A(n9536), .S(N22), .Y(n10487) );
  MUX2X1 U12641 ( .B(\RF[30][34] ), .A(\RF[31][34] ), .S(n10584), .Y(n9556) );
  MUX2X1 U12642 ( .B(\RF[28][34] ), .A(\RF[29][34] ), .S(n10584), .Y(n9555) );
  MUX2X1 U12643 ( .B(\RF[26][34] ), .A(\RF[27][34] ), .S(n10584), .Y(n9559) );
  MUX2X1 U12644 ( .B(\RF[24][34] ), .A(\RF[25][34] ), .S(n10584), .Y(n9558) );
  MUX2X1 U12645 ( .B(n9557), .A(n9554), .S(n10694), .Y(n9568) );
  MUX2X1 U12646 ( .B(\RF[22][34] ), .A(\RF[23][34] ), .S(n10584), .Y(n9562) );
  MUX2X1 U12647 ( .B(\RF[20][34] ), .A(\RF[21][34] ), .S(n10584), .Y(n9561) );
  MUX2X1 U12648 ( .B(\RF[18][34] ), .A(\RF[19][34] ), .S(n10584), .Y(n9565) );
  MUX2X1 U12649 ( .B(\RF[16][34] ), .A(\RF[17][34] ), .S(n10584), .Y(n9564) );
  MUX2X1 U12650 ( .B(n9563), .A(n9560), .S(n10694), .Y(n9567) );
  MUX2X1 U12651 ( .B(\RF[14][34] ), .A(\RF[15][34] ), .S(n10584), .Y(n9571) );
  MUX2X1 U12652 ( .B(\RF[12][34] ), .A(\RF[13][34] ), .S(n10584), .Y(n9570) );
  MUX2X1 U12653 ( .B(\RF[10][34] ), .A(\RF[11][34] ), .S(n10584), .Y(n9574) );
  MUX2X1 U12654 ( .B(\RF[8][34] ), .A(\RF[9][34] ), .S(n10584), .Y(n9573) );
  MUX2X1 U12655 ( .B(n9572), .A(n9569), .S(n10694), .Y(n9583) );
  MUX2X1 U12656 ( .B(\RF[6][34] ), .A(\RF[7][34] ), .S(n10585), .Y(n9577) );
  MUX2X1 U12657 ( .B(\RF[4][34] ), .A(\RF[5][34] ), .S(n10585), .Y(n9576) );
  MUX2X1 U12658 ( .B(\RF[2][34] ), .A(\RF[3][34] ), .S(n10585), .Y(n9580) );
  MUX2X1 U12659 ( .B(\RF[0][34] ), .A(\RF[1][34] ), .S(n10585), .Y(n9579) );
  MUX2X1 U12660 ( .B(n9578), .A(n9575), .S(n10694), .Y(n9582) );
  MUX2X1 U12661 ( .B(n9581), .A(n9566), .S(N22), .Y(n10488) );
  MUX2X1 U12662 ( .B(\RF[30][35] ), .A(\RF[31][35] ), .S(n10585), .Y(n9586) );
  MUX2X1 U12663 ( .B(\RF[28][35] ), .A(\RF[29][35] ), .S(n10585), .Y(n9585) );
  MUX2X1 U12664 ( .B(\RF[26][35] ), .A(\RF[27][35] ), .S(n10585), .Y(n9589) );
  MUX2X1 U12665 ( .B(\RF[24][35] ), .A(\RF[25][35] ), .S(n10585), .Y(n9588) );
  MUX2X1 U12666 ( .B(n9587), .A(n9584), .S(n10694), .Y(n9598) );
  MUX2X1 U12667 ( .B(\RF[22][35] ), .A(\RF[23][35] ), .S(n10585), .Y(n9592) );
  MUX2X1 U12668 ( .B(\RF[20][35] ), .A(\RF[21][35] ), .S(n10585), .Y(n9591) );
  MUX2X1 U12669 ( .B(\RF[18][35] ), .A(\RF[19][35] ), .S(n10585), .Y(n9595) );
  MUX2X1 U12670 ( .B(\RF[16][35] ), .A(\RF[17][35] ), .S(n10585), .Y(n9594) );
  MUX2X1 U12671 ( .B(n9593), .A(n9590), .S(n10694), .Y(n9597) );
  MUX2X1 U12672 ( .B(\RF[14][35] ), .A(\RF[15][35] ), .S(n10586), .Y(n9601) );
  MUX2X1 U12673 ( .B(\RF[12][35] ), .A(\RF[13][35] ), .S(n10586), .Y(n9600) );
  MUX2X1 U12674 ( .B(\RF[10][35] ), .A(\RF[11][35] ), .S(n10586), .Y(n9604) );
  MUX2X1 U12675 ( .B(\RF[8][35] ), .A(\RF[9][35] ), .S(n10586), .Y(n9603) );
  MUX2X1 U12676 ( .B(n9602), .A(n9599), .S(n10694), .Y(n9613) );
  MUX2X1 U12677 ( .B(\RF[6][35] ), .A(\RF[7][35] ), .S(n10586), .Y(n9607) );
  MUX2X1 U12678 ( .B(\RF[4][35] ), .A(\RF[5][35] ), .S(n10586), .Y(n9606) );
  MUX2X1 U12679 ( .B(\RF[2][35] ), .A(\RF[3][35] ), .S(n10586), .Y(n9610) );
  MUX2X1 U12680 ( .B(\RF[0][35] ), .A(\RF[1][35] ), .S(n10586), .Y(n9609) );
  MUX2X1 U12681 ( .B(n9608), .A(n9605), .S(n10694), .Y(n9612) );
  MUX2X1 U12682 ( .B(n9611), .A(n9596), .S(N22), .Y(n10489) );
  MUX2X1 U12683 ( .B(\RF[30][36] ), .A(\RF[31][36] ), .S(n10586), .Y(n9616) );
  MUX2X1 U12684 ( .B(\RF[28][36] ), .A(\RF[29][36] ), .S(n10586), .Y(n9615) );
  MUX2X1 U12685 ( .B(\RF[26][36] ), .A(\RF[27][36] ), .S(n10586), .Y(n9619) );
  MUX2X1 U12686 ( .B(\RF[24][36] ), .A(\RF[25][36] ), .S(n10586), .Y(n9618) );
  MUX2X1 U12687 ( .B(n9617), .A(n9614), .S(n10694), .Y(n9628) );
  MUX2X1 U12688 ( .B(\RF[22][36] ), .A(\RF[23][36] ), .S(n10587), .Y(n9622) );
  MUX2X1 U12689 ( .B(\RF[20][36] ), .A(\RF[21][36] ), .S(n10587), .Y(n9621) );
  MUX2X1 U12690 ( .B(\RF[18][36] ), .A(\RF[19][36] ), .S(n10587), .Y(n9625) );
  MUX2X1 U12691 ( .B(\RF[16][36] ), .A(\RF[17][36] ), .S(n10587), .Y(n9624) );
  MUX2X1 U12692 ( .B(n9623), .A(n9620), .S(n10694), .Y(n9627) );
  MUX2X1 U12693 ( .B(\RF[14][36] ), .A(\RF[15][36] ), .S(n10587), .Y(n9631) );
  MUX2X1 U12694 ( .B(\RF[12][36] ), .A(\RF[13][36] ), .S(n10587), .Y(n9630) );
  MUX2X1 U12695 ( .B(\RF[10][36] ), .A(\RF[11][36] ), .S(n10587), .Y(n9634) );
  MUX2X1 U12696 ( .B(\RF[8][36] ), .A(\RF[9][36] ), .S(n10587), .Y(n9633) );
  MUX2X1 U12697 ( .B(n9632), .A(n9629), .S(n10694), .Y(n9643) );
  MUX2X1 U12698 ( .B(\RF[6][36] ), .A(\RF[7][36] ), .S(n10587), .Y(n9637) );
  MUX2X1 U12699 ( .B(\RF[4][36] ), .A(\RF[5][36] ), .S(n10587), .Y(n9636) );
  MUX2X1 U12700 ( .B(\RF[2][36] ), .A(\RF[3][36] ), .S(n10587), .Y(n9640) );
  MUX2X1 U12701 ( .B(\RF[0][36] ), .A(\RF[1][36] ), .S(n10587), .Y(n9639) );
  MUX2X1 U12702 ( .B(n9638), .A(n9635), .S(n10694), .Y(n9642) );
  MUX2X1 U12703 ( .B(n9641), .A(n9626), .S(N22), .Y(n10490) );
  MUX2X1 U12704 ( .B(\RF[30][37] ), .A(\RF[31][37] ), .S(n10588), .Y(n9646) );
  MUX2X1 U12705 ( .B(\RF[28][37] ), .A(\RF[29][37] ), .S(n10588), .Y(n9645) );
  MUX2X1 U12706 ( .B(\RF[26][37] ), .A(\RF[27][37] ), .S(n10588), .Y(n9649) );
  MUX2X1 U12707 ( .B(\RF[24][37] ), .A(\RF[25][37] ), .S(n10588), .Y(n9648) );
  MUX2X1 U12708 ( .B(n9647), .A(n9644), .S(n10695), .Y(n9658) );
  MUX2X1 U12709 ( .B(\RF[22][37] ), .A(\RF[23][37] ), .S(n10588), .Y(n9652) );
  MUX2X1 U12710 ( .B(\RF[20][37] ), .A(\RF[21][37] ), .S(n10588), .Y(n9651) );
  MUX2X1 U12711 ( .B(\RF[18][37] ), .A(\RF[19][37] ), .S(n10588), .Y(n9655) );
  MUX2X1 U12712 ( .B(\RF[16][37] ), .A(\RF[17][37] ), .S(n10588), .Y(n9654) );
  MUX2X1 U12713 ( .B(n9653), .A(n9650), .S(n10695), .Y(n9657) );
  MUX2X1 U12714 ( .B(\RF[14][37] ), .A(\RF[15][37] ), .S(n10588), .Y(n9661) );
  MUX2X1 U12715 ( .B(\RF[12][37] ), .A(\RF[13][37] ), .S(n10588), .Y(n9660) );
  MUX2X1 U12716 ( .B(\RF[10][37] ), .A(\RF[11][37] ), .S(n10588), .Y(n9664) );
  MUX2X1 U12717 ( .B(\RF[8][37] ), .A(\RF[9][37] ), .S(n10588), .Y(n9663) );
  MUX2X1 U12718 ( .B(n9662), .A(n9659), .S(n10695), .Y(n9673) );
  MUX2X1 U12719 ( .B(\RF[6][37] ), .A(\RF[7][37] ), .S(n10589), .Y(n9667) );
  MUX2X1 U12720 ( .B(\RF[4][37] ), .A(\RF[5][37] ), .S(n10589), .Y(n9666) );
  MUX2X1 U12721 ( .B(\RF[2][37] ), .A(\RF[3][37] ), .S(n10589), .Y(n9670) );
  MUX2X1 U12722 ( .B(\RF[0][37] ), .A(\RF[1][37] ), .S(n10589), .Y(n9669) );
  MUX2X1 U12723 ( .B(n9668), .A(n9665), .S(n10695), .Y(n9672) );
  MUX2X1 U12724 ( .B(n9671), .A(n9656), .S(N22), .Y(n10491) );
  MUX2X1 U12725 ( .B(\RF[30][38] ), .A(\RF[31][38] ), .S(n10589), .Y(n9676) );
  MUX2X1 U12726 ( .B(\RF[28][38] ), .A(\RF[29][38] ), .S(n10589), .Y(n9675) );
  MUX2X1 U12727 ( .B(\RF[26][38] ), .A(\RF[27][38] ), .S(n10589), .Y(n9679) );
  MUX2X1 U12728 ( .B(\RF[24][38] ), .A(\RF[25][38] ), .S(n10589), .Y(n9678) );
  MUX2X1 U12729 ( .B(n9677), .A(n9674), .S(n10695), .Y(n9688) );
  MUX2X1 U12730 ( .B(\RF[22][38] ), .A(\RF[23][38] ), .S(n10589), .Y(n9682) );
  MUX2X1 U12731 ( .B(\RF[20][38] ), .A(\RF[21][38] ), .S(n10589), .Y(n9681) );
  MUX2X1 U12732 ( .B(\RF[18][38] ), .A(\RF[19][38] ), .S(n10589), .Y(n9685) );
  MUX2X1 U12733 ( .B(\RF[16][38] ), .A(\RF[17][38] ), .S(n10589), .Y(n9684) );
  MUX2X1 U12734 ( .B(n9683), .A(n9680), .S(n10695), .Y(n9687) );
  MUX2X1 U12735 ( .B(\RF[14][38] ), .A(\RF[15][38] ), .S(n10590), .Y(n9691) );
  MUX2X1 U12736 ( .B(\RF[12][38] ), .A(\RF[13][38] ), .S(n10590), .Y(n9690) );
  MUX2X1 U12737 ( .B(\RF[10][38] ), .A(\RF[11][38] ), .S(n10590), .Y(n9694) );
  MUX2X1 U12738 ( .B(\RF[8][38] ), .A(\RF[9][38] ), .S(n10590), .Y(n9693) );
  MUX2X1 U12739 ( .B(n9692), .A(n9689), .S(n10695), .Y(n9703) );
  MUX2X1 U12740 ( .B(\RF[6][38] ), .A(\RF[7][38] ), .S(n10590), .Y(n9697) );
  MUX2X1 U12741 ( .B(\RF[4][38] ), .A(\RF[5][38] ), .S(n10590), .Y(n9696) );
  MUX2X1 U12742 ( .B(\RF[2][38] ), .A(\RF[3][38] ), .S(n10590), .Y(n9700) );
  MUX2X1 U12743 ( .B(\RF[0][38] ), .A(\RF[1][38] ), .S(n10590), .Y(n9699) );
  MUX2X1 U12744 ( .B(n9698), .A(n9695), .S(n10695), .Y(n9702) );
  MUX2X1 U12745 ( .B(n9701), .A(n9686), .S(N22), .Y(n10492) );
  MUX2X1 U12746 ( .B(\RF[30][39] ), .A(\RF[31][39] ), .S(n10590), .Y(n9706) );
  MUX2X1 U12747 ( .B(\RF[28][39] ), .A(\RF[29][39] ), .S(n10590), .Y(n9705) );
  MUX2X1 U12748 ( .B(\RF[26][39] ), .A(\RF[27][39] ), .S(n10590), .Y(n9709) );
  MUX2X1 U12749 ( .B(\RF[24][39] ), .A(\RF[25][39] ), .S(n10590), .Y(n9708) );
  MUX2X1 U12750 ( .B(n9707), .A(n9704), .S(n10695), .Y(n9718) );
  MUX2X1 U12751 ( .B(\RF[22][39] ), .A(\RF[23][39] ), .S(n10591), .Y(n9712) );
  MUX2X1 U12752 ( .B(\RF[20][39] ), .A(\RF[21][39] ), .S(n10591), .Y(n9711) );
  MUX2X1 U12753 ( .B(\RF[18][39] ), .A(\RF[19][39] ), .S(n10591), .Y(n9715) );
  MUX2X1 U12754 ( .B(\RF[16][39] ), .A(\RF[17][39] ), .S(n10591), .Y(n9714) );
  MUX2X1 U12755 ( .B(n9713), .A(n9710), .S(n10695), .Y(n9717) );
  MUX2X1 U12756 ( .B(\RF[14][39] ), .A(\RF[15][39] ), .S(n10591), .Y(n9721) );
  MUX2X1 U12757 ( .B(\RF[12][39] ), .A(\RF[13][39] ), .S(n10591), .Y(n9720) );
  MUX2X1 U12758 ( .B(\RF[10][39] ), .A(\RF[11][39] ), .S(n10591), .Y(n9724) );
  MUX2X1 U12759 ( .B(\RF[8][39] ), .A(\RF[9][39] ), .S(n10591), .Y(n9723) );
  MUX2X1 U12760 ( .B(n9722), .A(n9719), .S(n10695), .Y(n9733) );
  MUX2X1 U12761 ( .B(\RF[6][39] ), .A(\RF[7][39] ), .S(n10591), .Y(n9727) );
  MUX2X1 U12762 ( .B(\RF[4][39] ), .A(\RF[5][39] ), .S(n10591), .Y(n9726) );
  MUX2X1 U12763 ( .B(\RF[2][39] ), .A(\RF[3][39] ), .S(n10591), .Y(n9730) );
  MUX2X1 U12764 ( .B(\RF[0][39] ), .A(\RF[1][39] ), .S(n10591), .Y(n9729) );
  MUX2X1 U12765 ( .B(n9728), .A(n9725), .S(n10695), .Y(n9732) );
  MUX2X1 U12766 ( .B(n9731), .A(n9716), .S(N22), .Y(n10493) );
  MUX2X1 U12767 ( .B(\RF[30][40] ), .A(\RF[31][40] ), .S(n10592), .Y(n9736) );
  MUX2X1 U12768 ( .B(\RF[28][40] ), .A(\RF[29][40] ), .S(n10592), .Y(n9735) );
  MUX2X1 U12769 ( .B(\RF[26][40] ), .A(\RF[27][40] ), .S(n10592), .Y(n9739) );
  MUX2X1 U12770 ( .B(\RF[24][40] ), .A(\RF[25][40] ), .S(n10592), .Y(n9738) );
  MUX2X1 U12771 ( .B(n9737), .A(n9734), .S(n10696), .Y(n9748) );
  MUX2X1 U12772 ( .B(\RF[22][40] ), .A(\RF[23][40] ), .S(n10592), .Y(n9742) );
  MUX2X1 U12773 ( .B(\RF[20][40] ), .A(\RF[21][40] ), .S(n10592), .Y(n9741) );
  MUX2X1 U12774 ( .B(\RF[18][40] ), .A(\RF[19][40] ), .S(n10592), .Y(n9745) );
  MUX2X1 U12775 ( .B(\RF[16][40] ), .A(\RF[17][40] ), .S(n10592), .Y(n9744) );
  MUX2X1 U12776 ( .B(n9743), .A(n9740), .S(n10696), .Y(n9747) );
  MUX2X1 U12777 ( .B(\RF[14][40] ), .A(\RF[15][40] ), .S(n10592), .Y(n9751) );
  MUX2X1 U12778 ( .B(\RF[12][40] ), .A(\RF[13][40] ), .S(n10592), .Y(n9750) );
  MUX2X1 U12779 ( .B(\RF[10][40] ), .A(\RF[11][40] ), .S(n10592), .Y(n9754) );
  MUX2X1 U12780 ( .B(\RF[8][40] ), .A(\RF[9][40] ), .S(n10592), .Y(n9753) );
  MUX2X1 U12781 ( .B(n9752), .A(n9749), .S(n10696), .Y(n9763) );
  MUX2X1 U12782 ( .B(\RF[6][40] ), .A(\RF[7][40] ), .S(n10593), .Y(n9757) );
  MUX2X1 U12783 ( .B(\RF[4][40] ), .A(\RF[5][40] ), .S(n10593), .Y(n9756) );
  MUX2X1 U12784 ( .B(\RF[2][40] ), .A(\RF[3][40] ), .S(n10593), .Y(n9760) );
  MUX2X1 U12785 ( .B(\RF[0][40] ), .A(\RF[1][40] ), .S(n10593), .Y(n9759) );
  MUX2X1 U12786 ( .B(n9758), .A(n9755), .S(n10696), .Y(n9762) );
  MUX2X1 U12787 ( .B(n9761), .A(n9746), .S(N22), .Y(n10494) );
  MUX2X1 U12788 ( .B(\RF[30][41] ), .A(\RF[31][41] ), .S(n10593), .Y(n9766) );
  MUX2X1 U12789 ( .B(\RF[28][41] ), .A(\RF[29][41] ), .S(n10593), .Y(n9765) );
  MUX2X1 U12790 ( .B(\RF[26][41] ), .A(\RF[27][41] ), .S(n10593), .Y(n9769) );
  MUX2X1 U12791 ( .B(\RF[24][41] ), .A(\RF[25][41] ), .S(n10593), .Y(n9768) );
  MUX2X1 U12792 ( .B(n9767), .A(n9764), .S(n10696), .Y(n9778) );
  MUX2X1 U12793 ( .B(\RF[22][41] ), .A(\RF[23][41] ), .S(n10593), .Y(n9772) );
  MUX2X1 U12794 ( .B(\RF[20][41] ), .A(\RF[21][41] ), .S(n10593), .Y(n9771) );
  MUX2X1 U12795 ( .B(\RF[18][41] ), .A(\RF[19][41] ), .S(n10593), .Y(n9775) );
  MUX2X1 U12796 ( .B(\RF[16][41] ), .A(\RF[17][41] ), .S(n10593), .Y(n9774) );
  MUX2X1 U12797 ( .B(n9773), .A(n9770), .S(n10696), .Y(n9777) );
  MUX2X1 U12798 ( .B(\RF[14][41] ), .A(\RF[15][41] ), .S(n10594), .Y(n9781) );
  MUX2X1 U12799 ( .B(\RF[12][41] ), .A(\RF[13][41] ), .S(n10594), .Y(n9780) );
  MUX2X1 U12800 ( .B(\RF[10][41] ), .A(\RF[11][41] ), .S(n10594), .Y(n9784) );
  MUX2X1 U12801 ( .B(\RF[8][41] ), .A(\RF[9][41] ), .S(n10594), .Y(n9783) );
  MUX2X1 U12802 ( .B(n9782), .A(n9779), .S(n10696), .Y(n9793) );
  MUX2X1 U12803 ( .B(\RF[6][41] ), .A(\RF[7][41] ), .S(n10594), .Y(n9787) );
  MUX2X1 U12804 ( .B(\RF[4][41] ), .A(\RF[5][41] ), .S(n10594), .Y(n9786) );
  MUX2X1 U12805 ( .B(\RF[2][41] ), .A(\RF[3][41] ), .S(n10594), .Y(n9790) );
  MUX2X1 U12806 ( .B(\RF[0][41] ), .A(\RF[1][41] ), .S(n10594), .Y(n9789) );
  MUX2X1 U12807 ( .B(n9788), .A(n9785), .S(n10696), .Y(n9792) );
  MUX2X1 U12808 ( .B(n9791), .A(n9776), .S(N22), .Y(n10495) );
  MUX2X1 U12809 ( .B(\RF[30][42] ), .A(\RF[31][42] ), .S(n10594), .Y(n9796) );
  MUX2X1 U12810 ( .B(\RF[28][42] ), .A(\RF[29][42] ), .S(n10594), .Y(n9795) );
  MUX2X1 U12811 ( .B(\RF[26][42] ), .A(\RF[27][42] ), .S(n10594), .Y(n9799) );
  MUX2X1 U12812 ( .B(\RF[24][42] ), .A(\RF[25][42] ), .S(n10594), .Y(n9798) );
  MUX2X1 U12813 ( .B(n9797), .A(n9794), .S(n10696), .Y(n9808) );
  MUX2X1 U12814 ( .B(\RF[22][42] ), .A(\RF[23][42] ), .S(n10595), .Y(n9802) );
  MUX2X1 U12815 ( .B(\RF[20][42] ), .A(\RF[21][42] ), .S(n10595), .Y(n9801) );
  MUX2X1 U12816 ( .B(\RF[18][42] ), .A(\RF[19][42] ), .S(n10595), .Y(n9805) );
  MUX2X1 U12817 ( .B(\RF[16][42] ), .A(\RF[17][42] ), .S(n10595), .Y(n9804) );
  MUX2X1 U12818 ( .B(n9803), .A(n9800), .S(n10696), .Y(n9807) );
  MUX2X1 U12819 ( .B(\RF[14][42] ), .A(\RF[15][42] ), .S(n10595), .Y(n9811) );
  MUX2X1 U12820 ( .B(\RF[12][42] ), .A(\RF[13][42] ), .S(n10595), .Y(n9810) );
  MUX2X1 U12821 ( .B(\RF[10][42] ), .A(\RF[11][42] ), .S(n10595), .Y(n9814) );
  MUX2X1 U12822 ( .B(\RF[8][42] ), .A(\RF[9][42] ), .S(n10595), .Y(n9813) );
  MUX2X1 U12823 ( .B(n9812), .A(n9809), .S(n10696), .Y(n9823) );
  MUX2X1 U12824 ( .B(\RF[6][42] ), .A(\RF[7][42] ), .S(n10595), .Y(n9817) );
  MUX2X1 U12825 ( .B(\RF[4][42] ), .A(\RF[5][42] ), .S(n10595), .Y(n9816) );
  MUX2X1 U12826 ( .B(\RF[2][42] ), .A(\RF[3][42] ), .S(n10595), .Y(n9820) );
  MUX2X1 U12827 ( .B(\RF[0][42] ), .A(\RF[1][42] ), .S(n10595), .Y(n9819) );
  MUX2X1 U12828 ( .B(n9818), .A(n9815), .S(n10696), .Y(n9822) );
  MUX2X1 U12829 ( .B(n9821), .A(n9806), .S(N22), .Y(n10496) );
  MUX2X1 U12830 ( .B(\RF[30][43] ), .A(\RF[31][43] ), .S(n10596), .Y(n9826) );
  MUX2X1 U12831 ( .B(\RF[28][43] ), .A(\RF[29][43] ), .S(n10596), .Y(n9825) );
  MUX2X1 U12832 ( .B(\RF[26][43] ), .A(\RF[27][43] ), .S(n10596), .Y(n9829) );
  MUX2X1 U12833 ( .B(\RF[24][43] ), .A(\RF[25][43] ), .S(n10596), .Y(n9828) );
  MUX2X1 U12834 ( .B(n9827), .A(n9824), .S(n10697), .Y(n9838) );
  MUX2X1 U12835 ( .B(\RF[22][43] ), .A(\RF[23][43] ), .S(n10596), .Y(n9832) );
  MUX2X1 U12836 ( .B(\RF[20][43] ), .A(\RF[21][43] ), .S(n10596), .Y(n9831) );
  MUX2X1 U12837 ( .B(\RF[18][43] ), .A(\RF[19][43] ), .S(n10596), .Y(n9835) );
  MUX2X1 U12838 ( .B(\RF[16][43] ), .A(\RF[17][43] ), .S(n10596), .Y(n9834) );
  MUX2X1 U12839 ( .B(n9833), .A(n9830), .S(n10697), .Y(n9837) );
  MUX2X1 U12840 ( .B(\RF[14][43] ), .A(\RF[15][43] ), .S(n10596), .Y(n9841) );
  MUX2X1 U12841 ( .B(\RF[12][43] ), .A(\RF[13][43] ), .S(n10596), .Y(n9840) );
  MUX2X1 U12842 ( .B(\RF[10][43] ), .A(\RF[11][43] ), .S(n10596), .Y(n9844) );
  MUX2X1 U12843 ( .B(\RF[8][43] ), .A(\RF[9][43] ), .S(n10596), .Y(n9843) );
  MUX2X1 U12844 ( .B(n9842), .A(n9839), .S(n10697), .Y(n9853) );
  MUX2X1 U12845 ( .B(\RF[6][43] ), .A(\RF[7][43] ), .S(n10597), .Y(n9847) );
  MUX2X1 U12846 ( .B(\RF[4][43] ), .A(\RF[5][43] ), .S(n10597), .Y(n9846) );
  MUX2X1 U12847 ( .B(\RF[2][43] ), .A(\RF[3][43] ), .S(n10597), .Y(n9850) );
  MUX2X1 U12848 ( .B(\RF[0][43] ), .A(\RF[1][43] ), .S(n10597), .Y(n9849) );
  MUX2X1 U12849 ( .B(n9848), .A(n9845), .S(n10697), .Y(n9852) );
  MUX2X1 U12850 ( .B(n9851), .A(n9836), .S(N22), .Y(n10497) );
  MUX2X1 U12851 ( .B(\RF[30][44] ), .A(\RF[31][44] ), .S(n10597), .Y(n9856) );
  MUX2X1 U12852 ( .B(\RF[28][44] ), .A(\RF[29][44] ), .S(n10597), .Y(n9855) );
  MUX2X1 U12853 ( .B(\RF[26][44] ), .A(\RF[27][44] ), .S(n10597), .Y(n9859) );
  MUX2X1 U12854 ( .B(\RF[24][44] ), .A(\RF[25][44] ), .S(n10597), .Y(n9858) );
  MUX2X1 U12855 ( .B(n9857), .A(n9854), .S(n10697), .Y(n9868) );
  MUX2X1 U12856 ( .B(\RF[22][44] ), .A(\RF[23][44] ), .S(n10597), .Y(n9862) );
  MUX2X1 U12857 ( .B(\RF[20][44] ), .A(\RF[21][44] ), .S(n10597), .Y(n9861) );
  MUX2X1 U12858 ( .B(\RF[18][44] ), .A(\RF[19][44] ), .S(n10597), .Y(n9865) );
  MUX2X1 U12859 ( .B(\RF[16][44] ), .A(\RF[17][44] ), .S(n10597), .Y(n9864) );
  MUX2X1 U12860 ( .B(n9863), .A(n9860), .S(n10697), .Y(n9867) );
  MUX2X1 U12861 ( .B(\RF[14][44] ), .A(\RF[15][44] ), .S(n10598), .Y(n9871) );
  MUX2X1 U12862 ( .B(\RF[12][44] ), .A(\RF[13][44] ), .S(n10598), .Y(n9870) );
  MUX2X1 U12863 ( .B(\RF[10][44] ), .A(\RF[11][44] ), .S(n10598), .Y(n9874) );
  MUX2X1 U12864 ( .B(\RF[8][44] ), .A(\RF[9][44] ), .S(n10598), .Y(n9873) );
  MUX2X1 U12865 ( .B(n9872), .A(n9869), .S(n10697), .Y(n9883) );
  MUX2X1 U12866 ( .B(\RF[6][44] ), .A(\RF[7][44] ), .S(n10598), .Y(n9877) );
  MUX2X1 U12867 ( .B(\RF[4][44] ), .A(\RF[5][44] ), .S(n10598), .Y(n9876) );
  MUX2X1 U12868 ( .B(\RF[2][44] ), .A(\RF[3][44] ), .S(n10598), .Y(n9880) );
  MUX2X1 U12869 ( .B(\RF[0][44] ), .A(\RF[1][44] ), .S(n10598), .Y(n9879) );
  MUX2X1 U12870 ( .B(n9878), .A(n9875), .S(n10697), .Y(n9882) );
  MUX2X1 U12871 ( .B(n9881), .A(n9866), .S(N22), .Y(n10498) );
  MUX2X1 U12872 ( .B(\RF[30][45] ), .A(\RF[31][45] ), .S(n10598), .Y(n9886) );
  MUX2X1 U12873 ( .B(\RF[28][45] ), .A(\RF[29][45] ), .S(n10598), .Y(n9885) );
  MUX2X1 U12874 ( .B(\RF[26][45] ), .A(\RF[27][45] ), .S(n10598), .Y(n9889) );
  MUX2X1 U12875 ( .B(\RF[24][45] ), .A(\RF[25][45] ), .S(n10598), .Y(n9888) );
  MUX2X1 U12876 ( .B(n9887), .A(n9884), .S(n10697), .Y(n9898) );
  MUX2X1 U12877 ( .B(\RF[22][45] ), .A(\RF[23][45] ), .S(n10599), .Y(n9892) );
  MUX2X1 U12878 ( .B(\RF[20][45] ), .A(\RF[21][45] ), .S(n10599), .Y(n9891) );
  MUX2X1 U12879 ( .B(\RF[18][45] ), .A(\RF[19][45] ), .S(n10599), .Y(n9895) );
  MUX2X1 U12880 ( .B(\RF[16][45] ), .A(\RF[17][45] ), .S(n10599), .Y(n9894) );
  MUX2X1 U12881 ( .B(n9893), .A(n9890), .S(n10697), .Y(n9897) );
  MUX2X1 U12882 ( .B(\RF[14][45] ), .A(\RF[15][45] ), .S(n10599), .Y(n9901) );
  MUX2X1 U12883 ( .B(\RF[12][45] ), .A(\RF[13][45] ), .S(n10599), .Y(n9900) );
  MUX2X1 U12884 ( .B(\RF[10][45] ), .A(\RF[11][45] ), .S(n10599), .Y(n9904) );
  MUX2X1 U12885 ( .B(\RF[8][45] ), .A(\RF[9][45] ), .S(n10599), .Y(n9903) );
  MUX2X1 U12886 ( .B(n9902), .A(n9899), .S(n10697), .Y(n9913) );
  MUX2X1 U12887 ( .B(\RF[6][45] ), .A(\RF[7][45] ), .S(n10599), .Y(n9907) );
  MUX2X1 U12888 ( .B(\RF[4][45] ), .A(\RF[5][45] ), .S(n10599), .Y(n9906) );
  MUX2X1 U12889 ( .B(\RF[2][45] ), .A(\RF[3][45] ), .S(n10599), .Y(n9910) );
  MUX2X1 U12890 ( .B(\RF[0][45] ), .A(\RF[1][45] ), .S(n10599), .Y(n9909) );
  MUX2X1 U12891 ( .B(n9908), .A(n9905), .S(n10697), .Y(n9912) );
  MUX2X1 U12892 ( .B(n9911), .A(n9896), .S(N22), .Y(n10499) );
  MUX2X1 U12893 ( .B(\RF[30][46] ), .A(\RF[31][46] ), .S(n10600), .Y(n9916) );
  MUX2X1 U12894 ( .B(\RF[28][46] ), .A(\RF[29][46] ), .S(n10600), .Y(n9915) );
  MUX2X1 U12895 ( .B(\RF[26][46] ), .A(\RF[27][46] ), .S(n10600), .Y(n9919) );
  MUX2X1 U12896 ( .B(\RF[24][46] ), .A(\RF[25][46] ), .S(n10600), .Y(n9918) );
  MUX2X1 U12897 ( .B(n9917), .A(n9914), .S(n10698), .Y(n9928) );
  MUX2X1 U12898 ( .B(\RF[22][46] ), .A(\RF[23][46] ), .S(n10600), .Y(n9922) );
  MUX2X1 U12899 ( .B(\RF[20][46] ), .A(\RF[21][46] ), .S(n10600), .Y(n9921) );
  MUX2X1 U12900 ( .B(\RF[18][46] ), .A(\RF[19][46] ), .S(n10600), .Y(n9925) );
  MUX2X1 U12901 ( .B(\RF[16][46] ), .A(\RF[17][46] ), .S(n10600), .Y(n9924) );
  MUX2X1 U12902 ( .B(n9923), .A(n9920), .S(n10698), .Y(n9927) );
  MUX2X1 U12903 ( .B(\RF[14][46] ), .A(\RF[15][46] ), .S(n10600), .Y(n9931) );
  MUX2X1 U12904 ( .B(\RF[12][46] ), .A(\RF[13][46] ), .S(n10600), .Y(n9930) );
  MUX2X1 U12905 ( .B(\RF[10][46] ), .A(\RF[11][46] ), .S(n10600), .Y(n9934) );
  MUX2X1 U12906 ( .B(\RF[8][46] ), .A(\RF[9][46] ), .S(n10600), .Y(n9933) );
  MUX2X1 U12907 ( .B(n9932), .A(n9929), .S(n10698), .Y(n9943) );
  MUX2X1 U12908 ( .B(\RF[6][46] ), .A(\RF[7][46] ), .S(n10601), .Y(n9937) );
  MUX2X1 U12909 ( .B(\RF[4][46] ), .A(\RF[5][46] ), .S(n10601), .Y(n9936) );
  MUX2X1 U12910 ( .B(\RF[2][46] ), .A(\RF[3][46] ), .S(n10601), .Y(n9940) );
  MUX2X1 U12911 ( .B(\RF[0][46] ), .A(\RF[1][46] ), .S(n10601), .Y(n9939) );
  MUX2X1 U12912 ( .B(n9938), .A(n9935), .S(n10698), .Y(n9942) );
  MUX2X1 U12913 ( .B(n9941), .A(n9926), .S(N22), .Y(n10500) );
  MUX2X1 U12914 ( .B(\RF[30][47] ), .A(\RF[31][47] ), .S(n10601), .Y(n9946) );
  MUX2X1 U12915 ( .B(\RF[28][47] ), .A(\RF[29][47] ), .S(n10601), .Y(n9945) );
  MUX2X1 U12916 ( .B(\RF[26][47] ), .A(\RF[27][47] ), .S(n10601), .Y(n9949) );
  MUX2X1 U12917 ( .B(\RF[24][47] ), .A(\RF[25][47] ), .S(n10601), .Y(n9948) );
  MUX2X1 U12918 ( .B(n9947), .A(n9944), .S(n10698), .Y(n9958) );
  MUX2X1 U12919 ( .B(\RF[22][47] ), .A(\RF[23][47] ), .S(n10601), .Y(n9952) );
  MUX2X1 U12920 ( .B(\RF[20][47] ), .A(\RF[21][47] ), .S(n10601), .Y(n9951) );
  MUX2X1 U12921 ( .B(\RF[18][47] ), .A(\RF[19][47] ), .S(n10601), .Y(n9955) );
  MUX2X1 U12922 ( .B(\RF[16][47] ), .A(\RF[17][47] ), .S(n10601), .Y(n9954) );
  MUX2X1 U12923 ( .B(n9953), .A(n9950), .S(n10698), .Y(n9957) );
  MUX2X1 U12924 ( .B(\RF[14][47] ), .A(\RF[15][47] ), .S(n10602), .Y(n9961) );
  MUX2X1 U12925 ( .B(\RF[12][47] ), .A(\RF[13][47] ), .S(n10602), .Y(n9960) );
  MUX2X1 U12926 ( .B(\RF[10][47] ), .A(\RF[11][47] ), .S(n10602), .Y(n9964) );
  MUX2X1 U12927 ( .B(\RF[8][47] ), .A(\RF[9][47] ), .S(n10602), .Y(n9963) );
  MUX2X1 U12928 ( .B(n9962), .A(n9959), .S(n10698), .Y(n9973) );
  MUX2X1 U12929 ( .B(\RF[6][47] ), .A(\RF[7][47] ), .S(n10602), .Y(n9967) );
  MUX2X1 U12930 ( .B(\RF[4][47] ), .A(\RF[5][47] ), .S(n10602), .Y(n9966) );
  MUX2X1 U12931 ( .B(\RF[2][47] ), .A(\RF[3][47] ), .S(n10602), .Y(n9970) );
  MUX2X1 U12932 ( .B(\RF[0][47] ), .A(\RF[1][47] ), .S(n10602), .Y(n9969) );
  MUX2X1 U12933 ( .B(n9968), .A(n9965), .S(n10698), .Y(n9972) );
  MUX2X1 U12934 ( .B(n9971), .A(n9956), .S(N22), .Y(n10501) );
  MUX2X1 U12935 ( .B(\RF[30][48] ), .A(\RF[31][48] ), .S(n10602), .Y(n9976) );
  MUX2X1 U12936 ( .B(\RF[28][48] ), .A(\RF[29][48] ), .S(n10602), .Y(n9975) );
  MUX2X1 U12937 ( .B(\RF[26][48] ), .A(\RF[27][48] ), .S(n10602), .Y(n9979) );
  MUX2X1 U12938 ( .B(\RF[24][48] ), .A(\RF[25][48] ), .S(n10602), .Y(n9978) );
  MUX2X1 U12939 ( .B(n9977), .A(n9974), .S(n10698), .Y(n9988) );
  MUX2X1 U12940 ( .B(\RF[22][48] ), .A(\RF[23][48] ), .S(n10603), .Y(n9982) );
  MUX2X1 U12941 ( .B(\RF[20][48] ), .A(\RF[21][48] ), .S(n10603), .Y(n9981) );
  MUX2X1 U12942 ( .B(\RF[18][48] ), .A(\RF[19][48] ), .S(n10603), .Y(n9985) );
  MUX2X1 U12943 ( .B(\RF[16][48] ), .A(\RF[17][48] ), .S(n10603), .Y(n9984) );
  MUX2X1 U12944 ( .B(n9983), .A(n9980), .S(n10698), .Y(n9987) );
  MUX2X1 U12945 ( .B(\RF[14][48] ), .A(\RF[15][48] ), .S(n10603), .Y(n9991) );
  MUX2X1 U12946 ( .B(\RF[12][48] ), .A(\RF[13][48] ), .S(n10603), .Y(n9990) );
  MUX2X1 U12947 ( .B(\RF[10][48] ), .A(\RF[11][48] ), .S(n10603), .Y(n9994) );
  MUX2X1 U12948 ( .B(\RF[8][48] ), .A(\RF[9][48] ), .S(n10603), .Y(n9993) );
  MUX2X1 U12949 ( .B(n9992), .A(n9989), .S(n10698), .Y(n10003) );
  MUX2X1 U12950 ( .B(\RF[6][48] ), .A(\RF[7][48] ), .S(n10603), .Y(n9997) );
  MUX2X1 U12951 ( .B(\RF[4][48] ), .A(\RF[5][48] ), .S(n10603), .Y(n9996) );
  MUX2X1 U12952 ( .B(\RF[2][48] ), .A(\RF[3][48] ), .S(n10603), .Y(n10000) );
  MUX2X1 U12953 ( .B(\RF[0][48] ), .A(\RF[1][48] ), .S(n10603), .Y(n9999) );
  MUX2X1 U12954 ( .B(n9998), .A(n9995), .S(n10698), .Y(n10002) );
  MUX2X1 U12955 ( .B(n10001), .A(n9986), .S(N22), .Y(n10502) );
  MUX2X1 U12956 ( .B(\RF[30][49] ), .A(\RF[31][49] ), .S(n10604), .Y(n10006)
         );
  MUX2X1 U12957 ( .B(\RF[28][49] ), .A(\RF[29][49] ), .S(n10604), .Y(n10005)
         );
  MUX2X1 U12958 ( .B(\RF[26][49] ), .A(\RF[27][49] ), .S(n10604), .Y(n10009)
         );
  MUX2X1 U12959 ( .B(\RF[24][49] ), .A(\RF[25][49] ), .S(n10604), .Y(n10008)
         );
  MUX2X1 U12960 ( .B(n10007), .A(n10004), .S(n10694), .Y(n10018) );
  MUX2X1 U12961 ( .B(\RF[22][49] ), .A(\RF[23][49] ), .S(n10604), .Y(n10012)
         );
  MUX2X1 U12962 ( .B(\RF[20][49] ), .A(\RF[21][49] ), .S(n10604), .Y(n10011)
         );
  MUX2X1 U12963 ( .B(\RF[18][49] ), .A(\RF[19][49] ), .S(n10604), .Y(n10015)
         );
  MUX2X1 U12964 ( .B(\RF[16][49] ), .A(\RF[17][49] ), .S(n10604), .Y(n10014)
         );
  MUX2X1 U12965 ( .B(n10013), .A(n10010), .S(n10688), .Y(n10017) );
  MUX2X1 U12966 ( .B(\RF[14][49] ), .A(\RF[15][49] ), .S(n10604), .Y(n10021)
         );
  MUX2X1 U12967 ( .B(\RF[12][49] ), .A(\RF[13][49] ), .S(n10604), .Y(n10020)
         );
  MUX2X1 U12968 ( .B(\RF[10][49] ), .A(\RF[11][49] ), .S(n10604), .Y(n10024)
         );
  MUX2X1 U12969 ( .B(\RF[8][49] ), .A(\RF[9][49] ), .S(n10604), .Y(n10023) );
  MUX2X1 U12970 ( .B(n10022), .A(n10019), .S(n10690), .Y(n10033) );
  MUX2X1 U12971 ( .B(\RF[6][49] ), .A(\RF[7][49] ), .S(n10605), .Y(n10027) );
  MUX2X1 U12972 ( .B(\RF[4][49] ), .A(\RF[5][49] ), .S(n10605), .Y(n10026) );
  MUX2X1 U12973 ( .B(\RF[2][49] ), .A(\RF[3][49] ), .S(n10605), .Y(n10030) );
  MUX2X1 U12974 ( .B(\RF[0][49] ), .A(\RF[1][49] ), .S(n10605), .Y(n10029) );
  MUX2X1 U12975 ( .B(n10028), .A(n10025), .S(n10691), .Y(n10032) );
  MUX2X1 U12976 ( .B(n10031), .A(n10016), .S(N22), .Y(n10503) );
  MUX2X1 U12977 ( .B(\RF[30][50] ), .A(\RF[31][50] ), .S(n10605), .Y(n10036)
         );
  MUX2X1 U12978 ( .B(\RF[28][50] ), .A(\RF[29][50] ), .S(n10605), .Y(n10035)
         );
  MUX2X1 U12979 ( .B(\RF[26][50] ), .A(\RF[27][50] ), .S(n10605), .Y(n10039)
         );
  MUX2X1 U12980 ( .B(\RF[24][50] ), .A(\RF[25][50] ), .S(n10605), .Y(n10038)
         );
  MUX2X1 U12981 ( .B(n10037), .A(n10034), .S(n10696), .Y(n10048) );
  MUX2X1 U12982 ( .B(\RF[22][50] ), .A(\RF[23][50] ), .S(n10605), .Y(n10042)
         );
  MUX2X1 U12983 ( .B(\RF[20][50] ), .A(\RF[21][50] ), .S(n10605), .Y(n10041)
         );
  MUX2X1 U12984 ( .B(\RF[18][50] ), .A(\RF[19][50] ), .S(n10605), .Y(n10045)
         );
  MUX2X1 U12985 ( .B(\RF[16][50] ), .A(\RF[17][50] ), .S(n10605), .Y(n10044)
         );
  MUX2X1 U12986 ( .B(n10043), .A(n10040), .S(n10686), .Y(n10047) );
  MUX2X1 U12987 ( .B(\RF[14][50] ), .A(\RF[15][50] ), .S(n10606), .Y(n10051)
         );
  MUX2X1 U12988 ( .B(\RF[12][50] ), .A(\RF[13][50] ), .S(n10606), .Y(n10050)
         );
  MUX2X1 U12989 ( .B(\RF[10][50] ), .A(\RF[11][50] ), .S(n10606), .Y(n10054)
         );
  MUX2X1 U12990 ( .B(\RF[8][50] ), .A(\RF[9][50] ), .S(n10606), .Y(n10053) );
  MUX2X1 U12991 ( .B(n10052), .A(n10049), .S(n10687), .Y(n10063) );
  MUX2X1 U12992 ( .B(\RF[6][50] ), .A(\RF[7][50] ), .S(n10606), .Y(n10057) );
  MUX2X1 U12993 ( .B(\RF[4][50] ), .A(\RF[5][50] ), .S(n10606), .Y(n10056) );
  MUX2X1 U12994 ( .B(\RF[2][50] ), .A(\RF[3][50] ), .S(n10606), .Y(n10060) );
  MUX2X1 U12995 ( .B(\RF[0][50] ), .A(\RF[1][50] ), .S(n10606), .Y(n10059) );
  MUX2X1 U12996 ( .B(n10058), .A(n10055), .S(N20), .Y(n10062) );
  MUX2X1 U12997 ( .B(n10061), .A(n10046), .S(N22), .Y(n10504) );
  MUX2X1 U12998 ( .B(\RF[30][51] ), .A(\RF[31][51] ), .S(n10606), .Y(n10066)
         );
  MUX2X1 U12999 ( .B(\RF[28][51] ), .A(\RF[29][51] ), .S(n10606), .Y(n10065)
         );
  MUX2X1 U13000 ( .B(\RF[26][51] ), .A(\RF[27][51] ), .S(n10606), .Y(n10069)
         );
  MUX2X1 U13001 ( .B(\RF[24][51] ), .A(\RF[25][51] ), .S(n10606), .Y(n10068)
         );
  MUX2X1 U13002 ( .B(n10067), .A(n10064), .S(n10692), .Y(n10078) );
  MUX2X1 U13003 ( .B(\RF[22][51] ), .A(\RF[23][51] ), .S(n10607), .Y(n10072)
         );
  MUX2X1 U13004 ( .B(\RF[20][51] ), .A(\RF[21][51] ), .S(n10607), .Y(n10071)
         );
  MUX2X1 U13005 ( .B(\RF[18][51] ), .A(\RF[19][51] ), .S(n10607), .Y(n10075)
         );
  MUX2X1 U13006 ( .B(\RF[16][51] ), .A(\RF[17][51] ), .S(n10607), .Y(n10074)
         );
  MUX2X1 U13007 ( .B(n10073), .A(n10070), .S(n10697), .Y(n10077) );
  MUX2X1 U13008 ( .B(\RF[14][51] ), .A(\RF[15][51] ), .S(n10607), .Y(n10081)
         );
  MUX2X1 U13009 ( .B(\RF[12][51] ), .A(\RF[13][51] ), .S(n10607), .Y(n10080)
         );
  MUX2X1 U13010 ( .B(\RF[10][51] ), .A(\RF[11][51] ), .S(n10607), .Y(n10084)
         );
  MUX2X1 U13011 ( .B(\RF[8][51] ), .A(\RF[9][51] ), .S(n10607), .Y(n10083) );
  MUX2X1 U13012 ( .B(n10082), .A(n10079), .S(n10689), .Y(n10093) );
  MUX2X1 U13013 ( .B(\RF[6][51] ), .A(\RF[7][51] ), .S(n10607), .Y(n10087) );
  MUX2X1 U13014 ( .B(\RF[4][51] ), .A(\RF[5][51] ), .S(n10607), .Y(n10086) );
  MUX2X1 U13015 ( .B(\RF[2][51] ), .A(\RF[3][51] ), .S(n10607), .Y(n10090) );
  MUX2X1 U13016 ( .B(\RF[0][51] ), .A(\RF[1][51] ), .S(n10607), .Y(n10089) );
  MUX2X1 U13017 ( .B(n10088), .A(n10085), .S(n10698), .Y(n10092) );
  MUX2X1 U13018 ( .B(n10091), .A(n10076), .S(N22), .Y(n10505) );
  MUX2X1 U13019 ( .B(\RF[30][52] ), .A(\RF[31][52] ), .S(n10608), .Y(n10096)
         );
  MUX2X1 U13020 ( .B(\RF[28][52] ), .A(\RF[29][52] ), .S(n10608), .Y(n10095)
         );
  MUX2X1 U13021 ( .B(\RF[26][52] ), .A(\RF[27][52] ), .S(n10608), .Y(n10099)
         );
  MUX2X1 U13022 ( .B(\RF[24][52] ), .A(\RF[25][52] ), .S(n10608), .Y(n10098)
         );
  MUX2X1 U13023 ( .B(n10097), .A(n10094), .S(n10699), .Y(n10108) );
  MUX2X1 U13024 ( .B(\RF[22][52] ), .A(\RF[23][52] ), .S(n10608), .Y(n10102)
         );
  MUX2X1 U13025 ( .B(\RF[20][52] ), .A(\RF[21][52] ), .S(n10608), .Y(n10101)
         );
  MUX2X1 U13026 ( .B(\RF[18][52] ), .A(\RF[19][52] ), .S(n10608), .Y(n10105)
         );
  MUX2X1 U13027 ( .B(\RF[16][52] ), .A(\RF[17][52] ), .S(n10608), .Y(n10104)
         );
  MUX2X1 U13028 ( .B(n10103), .A(n10100), .S(n10699), .Y(n10107) );
  MUX2X1 U13029 ( .B(\RF[14][52] ), .A(\RF[15][52] ), .S(n10608), .Y(n10111)
         );
  MUX2X1 U13030 ( .B(\RF[12][52] ), .A(\RF[13][52] ), .S(n10608), .Y(n10110)
         );
  MUX2X1 U13031 ( .B(\RF[10][52] ), .A(\RF[11][52] ), .S(n10608), .Y(n10114)
         );
  MUX2X1 U13032 ( .B(\RF[8][52] ), .A(\RF[9][52] ), .S(n10608), .Y(n10113) );
  MUX2X1 U13033 ( .B(n10112), .A(n10109), .S(n10699), .Y(n10123) );
  MUX2X1 U13034 ( .B(\RF[6][52] ), .A(\RF[7][52] ), .S(n10609), .Y(n10117) );
  MUX2X1 U13035 ( .B(\RF[4][52] ), .A(\RF[5][52] ), .S(n10609), .Y(n10116) );
  MUX2X1 U13036 ( .B(\RF[2][52] ), .A(\RF[3][52] ), .S(n10609), .Y(n10120) );
  MUX2X1 U13037 ( .B(\RF[0][52] ), .A(\RF[1][52] ), .S(n10609), .Y(n10119) );
  MUX2X1 U13038 ( .B(n10118), .A(n10115), .S(n10699), .Y(n10122) );
  MUX2X1 U13039 ( .B(n10121), .A(n10106), .S(N22), .Y(n10506) );
  MUX2X1 U13040 ( .B(\RF[30][53] ), .A(\RF[31][53] ), .S(n10609), .Y(n10126)
         );
  MUX2X1 U13041 ( .B(\RF[28][53] ), .A(\RF[29][53] ), .S(n10609), .Y(n10125)
         );
  MUX2X1 U13042 ( .B(\RF[26][53] ), .A(\RF[27][53] ), .S(n10609), .Y(n10129)
         );
  MUX2X1 U13043 ( .B(\RF[24][53] ), .A(\RF[25][53] ), .S(n10609), .Y(n10128)
         );
  MUX2X1 U13044 ( .B(n10127), .A(n10124), .S(n10699), .Y(n10138) );
  MUX2X1 U13045 ( .B(\RF[22][53] ), .A(\RF[23][53] ), .S(n10609), .Y(n10132)
         );
  MUX2X1 U13046 ( .B(\RF[20][53] ), .A(\RF[21][53] ), .S(n10609), .Y(n10131)
         );
  MUX2X1 U13047 ( .B(\RF[18][53] ), .A(\RF[19][53] ), .S(n10609), .Y(n10135)
         );
  MUX2X1 U13048 ( .B(\RF[16][53] ), .A(\RF[17][53] ), .S(n10609), .Y(n10134)
         );
  MUX2X1 U13049 ( .B(n10133), .A(n10130), .S(n10699), .Y(n10137) );
  MUX2X1 U13050 ( .B(\RF[14][53] ), .A(\RF[15][53] ), .S(n10610), .Y(n10141)
         );
  MUX2X1 U13051 ( .B(\RF[12][53] ), .A(\RF[13][53] ), .S(n10610), .Y(n10140)
         );
  MUX2X1 U13052 ( .B(\RF[10][53] ), .A(\RF[11][53] ), .S(n10610), .Y(n10144)
         );
  MUX2X1 U13053 ( .B(\RF[8][53] ), .A(\RF[9][53] ), .S(n10610), .Y(n10143) );
  MUX2X1 U13054 ( .B(n10142), .A(n10139), .S(n10699), .Y(n10153) );
  MUX2X1 U13055 ( .B(\RF[6][53] ), .A(\RF[7][53] ), .S(n10610), .Y(n10147) );
  MUX2X1 U13056 ( .B(\RF[4][53] ), .A(\RF[5][53] ), .S(n10610), .Y(n10146) );
  MUX2X1 U13057 ( .B(\RF[2][53] ), .A(\RF[3][53] ), .S(n10610), .Y(n10150) );
  MUX2X1 U13058 ( .B(\RF[0][53] ), .A(\RF[1][53] ), .S(n10610), .Y(n10149) );
  MUX2X1 U13059 ( .B(n10148), .A(n10145), .S(n10699), .Y(n10152) );
  MUX2X1 U13060 ( .B(n10151), .A(n10136), .S(N22), .Y(n10507) );
  MUX2X1 U13061 ( .B(\RF[30][54] ), .A(\RF[31][54] ), .S(n10610), .Y(n10156)
         );
  MUX2X1 U13062 ( .B(\RF[28][54] ), .A(\RF[29][54] ), .S(n10610), .Y(n10155)
         );
  MUX2X1 U13063 ( .B(\RF[26][54] ), .A(\RF[27][54] ), .S(n10610), .Y(n10159)
         );
  MUX2X1 U13064 ( .B(\RF[24][54] ), .A(\RF[25][54] ), .S(n10610), .Y(n10158)
         );
  MUX2X1 U13065 ( .B(n10157), .A(n10154), .S(n10699), .Y(n10168) );
  MUX2X1 U13066 ( .B(\RF[22][54] ), .A(\RF[23][54] ), .S(n10611), .Y(n10162)
         );
  MUX2X1 U13067 ( .B(\RF[20][54] ), .A(\RF[21][54] ), .S(n10611), .Y(n10161)
         );
  MUX2X1 U13068 ( .B(\RF[18][54] ), .A(\RF[19][54] ), .S(n10611), .Y(n10165)
         );
  MUX2X1 U13069 ( .B(\RF[16][54] ), .A(\RF[17][54] ), .S(n10611), .Y(n10164)
         );
  MUX2X1 U13070 ( .B(n10163), .A(n10160), .S(n10699), .Y(n10167) );
  MUX2X1 U13071 ( .B(\RF[14][54] ), .A(\RF[15][54] ), .S(n10611), .Y(n10171)
         );
  MUX2X1 U13072 ( .B(\RF[12][54] ), .A(\RF[13][54] ), .S(n10611), .Y(n10170)
         );
  MUX2X1 U13073 ( .B(\RF[10][54] ), .A(\RF[11][54] ), .S(n10611), .Y(n10174)
         );
  MUX2X1 U13074 ( .B(\RF[8][54] ), .A(\RF[9][54] ), .S(n10611), .Y(n10173) );
  MUX2X1 U13075 ( .B(n10172), .A(n10169), .S(n10699), .Y(n10183) );
  MUX2X1 U13076 ( .B(\RF[6][54] ), .A(\RF[7][54] ), .S(n10611), .Y(n10177) );
  MUX2X1 U13077 ( .B(\RF[4][54] ), .A(\RF[5][54] ), .S(n10611), .Y(n10176) );
  MUX2X1 U13078 ( .B(\RF[2][54] ), .A(\RF[3][54] ), .S(n10611), .Y(n10180) );
  MUX2X1 U13079 ( .B(\RF[0][54] ), .A(\RF[1][54] ), .S(n10611), .Y(n10179) );
  MUX2X1 U13080 ( .B(n10178), .A(n10175), .S(n10699), .Y(n10182) );
  MUX2X1 U13081 ( .B(n10181), .A(n10166), .S(N22), .Y(n10508) );
  MUX2X1 U13082 ( .B(\RF[30][55] ), .A(\RF[31][55] ), .S(n10612), .Y(n10186)
         );
  MUX2X1 U13083 ( .B(\RF[28][55] ), .A(\RF[29][55] ), .S(n10612), .Y(n10185)
         );
  MUX2X1 U13084 ( .B(\RF[26][55] ), .A(\RF[27][55] ), .S(n10612), .Y(n10189)
         );
  MUX2X1 U13085 ( .B(\RF[24][55] ), .A(\RF[25][55] ), .S(n10612), .Y(n10188)
         );
  MUX2X1 U13086 ( .B(n10187), .A(n10184), .S(n10700), .Y(n10198) );
  MUX2X1 U13087 ( .B(\RF[22][55] ), .A(\RF[23][55] ), .S(n10612), .Y(n10192)
         );
  MUX2X1 U13088 ( .B(\RF[20][55] ), .A(\RF[21][55] ), .S(n10612), .Y(n10191)
         );
  MUX2X1 U13089 ( .B(\RF[18][55] ), .A(\RF[19][55] ), .S(n10612), .Y(n10195)
         );
  MUX2X1 U13090 ( .B(\RF[16][55] ), .A(\RF[17][55] ), .S(n10612), .Y(n10194)
         );
  MUX2X1 U13091 ( .B(n10193), .A(n10190), .S(n10700), .Y(n10197) );
  MUX2X1 U13092 ( .B(\RF[14][55] ), .A(\RF[15][55] ), .S(n10612), .Y(n10201)
         );
  MUX2X1 U13093 ( .B(\RF[12][55] ), .A(\RF[13][55] ), .S(n10612), .Y(n10200)
         );
  MUX2X1 U13094 ( .B(\RF[10][55] ), .A(\RF[11][55] ), .S(n10612), .Y(n10204)
         );
  MUX2X1 U13095 ( .B(\RF[8][55] ), .A(\RF[9][55] ), .S(n10612), .Y(n10203) );
  MUX2X1 U13096 ( .B(n10202), .A(n10199), .S(n10700), .Y(n10213) );
  MUX2X1 U13097 ( .B(\RF[6][55] ), .A(\RF[7][55] ), .S(n10613), .Y(n10207) );
  MUX2X1 U13098 ( .B(\RF[4][55] ), .A(\RF[5][55] ), .S(n10613), .Y(n10206) );
  MUX2X1 U13099 ( .B(\RF[2][55] ), .A(\RF[3][55] ), .S(n10613), .Y(n10210) );
  MUX2X1 U13100 ( .B(\RF[0][55] ), .A(\RF[1][55] ), .S(n10613), .Y(n10209) );
  MUX2X1 U13101 ( .B(n10208), .A(n10205), .S(n10700), .Y(n10212) );
  MUX2X1 U13102 ( .B(n10211), .A(n10196), .S(N22), .Y(n10509) );
  MUX2X1 U13103 ( .B(\RF[30][56] ), .A(\RF[31][56] ), .S(n10613), .Y(n10216)
         );
  MUX2X1 U13104 ( .B(\RF[28][56] ), .A(\RF[29][56] ), .S(n10613), .Y(n10215)
         );
  MUX2X1 U13105 ( .B(\RF[26][56] ), .A(\RF[27][56] ), .S(n10613), .Y(n10219)
         );
  MUX2X1 U13106 ( .B(\RF[24][56] ), .A(\RF[25][56] ), .S(n10613), .Y(n10218)
         );
  MUX2X1 U13107 ( .B(n10217), .A(n10214), .S(n10700), .Y(n10228) );
  MUX2X1 U13108 ( .B(\RF[22][56] ), .A(\RF[23][56] ), .S(n10613), .Y(n10222)
         );
  MUX2X1 U13109 ( .B(\RF[20][56] ), .A(\RF[21][56] ), .S(n10613), .Y(n10221)
         );
  MUX2X1 U13110 ( .B(\RF[18][56] ), .A(\RF[19][56] ), .S(n10613), .Y(n10225)
         );
  MUX2X1 U13111 ( .B(\RF[16][56] ), .A(\RF[17][56] ), .S(n10613), .Y(n10224)
         );
  MUX2X1 U13112 ( .B(n10223), .A(n10220), .S(n10700), .Y(n10227) );
  MUX2X1 U13113 ( .B(\RF[14][56] ), .A(\RF[15][56] ), .S(n10614), .Y(n10231)
         );
  MUX2X1 U13114 ( .B(\RF[12][56] ), .A(\RF[13][56] ), .S(n10614), .Y(n10230)
         );
  MUX2X1 U13115 ( .B(\RF[10][56] ), .A(\RF[11][56] ), .S(n10614), .Y(n10234)
         );
  MUX2X1 U13116 ( .B(\RF[8][56] ), .A(\RF[9][56] ), .S(n10614), .Y(n10233) );
  MUX2X1 U13117 ( .B(n10232), .A(n10229), .S(n10700), .Y(n10243) );
  MUX2X1 U13118 ( .B(\RF[6][56] ), .A(\RF[7][56] ), .S(n10614), .Y(n10237) );
  MUX2X1 U13119 ( .B(\RF[4][56] ), .A(\RF[5][56] ), .S(n10614), .Y(n10236) );
  MUX2X1 U13120 ( .B(\RF[2][56] ), .A(\RF[3][56] ), .S(n10614), .Y(n10240) );
  MUX2X1 U13121 ( .B(\RF[0][56] ), .A(\RF[1][56] ), .S(n10614), .Y(n10239) );
  MUX2X1 U13122 ( .B(n10238), .A(n10235), .S(n10700), .Y(n10242) );
  MUX2X1 U13123 ( .B(n10241), .A(n10226), .S(N22), .Y(n10510) );
  MUX2X1 U13124 ( .B(\RF[30][57] ), .A(\RF[31][57] ), .S(n10614), .Y(n10246)
         );
  MUX2X1 U13125 ( .B(\RF[28][57] ), .A(\RF[29][57] ), .S(n10614), .Y(n10245)
         );
  MUX2X1 U13126 ( .B(\RF[26][57] ), .A(\RF[27][57] ), .S(n10614), .Y(n10249)
         );
  MUX2X1 U13127 ( .B(\RF[24][57] ), .A(\RF[25][57] ), .S(n10614), .Y(n10248)
         );
  MUX2X1 U13128 ( .B(n10247), .A(n10244), .S(n10700), .Y(n10258) );
  MUX2X1 U13129 ( .B(\RF[22][57] ), .A(\RF[23][57] ), .S(n10615), .Y(n10252)
         );
  MUX2X1 U13130 ( .B(\RF[20][57] ), .A(\RF[21][57] ), .S(n10615), .Y(n10251)
         );
  MUX2X1 U13131 ( .B(\RF[18][57] ), .A(\RF[19][57] ), .S(n10615), .Y(n10255)
         );
  MUX2X1 U13132 ( .B(\RF[16][57] ), .A(\RF[17][57] ), .S(n10615), .Y(n10254)
         );
  MUX2X1 U13133 ( .B(n10253), .A(n10250), .S(n10700), .Y(n10257) );
  MUX2X1 U13134 ( .B(\RF[14][57] ), .A(\RF[15][57] ), .S(n10615), .Y(n10261)
         );
  MUX2X1 U13135 ( .B(\RF[12][57] ), .A(\RF[13][57] ), .S(n10615), .Y(n10260)
         );
  MUX2X1 U13136 ( .B(\RF[10][57] ), .A(\RF[11][57] ), .S(n10615), .Y(n10264)
         );
  MUX2X1 U13137 ( .B(\RF[8][57] ), .A(\RF[9][57] ), .S(n10615), .Y(n10263) );
  MUX2X1 U13138 ( .B(n10262), .A(n10259), .S(n10700), .Y(n10273) );
  MUX2X1 U13139 ( .B(\RF[6][57] ), .A(\RF[7][57] ), .S(n10615), .Y(n10267) );
  MUX2X1 U13140 ( .B(\RF[4][57] ), .A(\RF[5][57] ), .S(n10615), .Y(n10266) );
  MUX2X1 U13141 ( .B(\RF[2][57] ), .A(\RF[3][57] ), .S(n10615), .Y(n10270) );
  MUX2X1 U13142 ( .B(\RF[0][57] ), .A(\RF[1][57] ), .S(n10615), .Y(n10269) );
  MUX2X1 U13143 ( .B(n10268), .A(n10265), .S(n10700), .Y(n10272) );
  MUX2X1 U13144 ( .B(n10271), .A(n10256), .S(N22), .Y(n10511) );
  MUX2X1 U13145 ( .B(\RF[30][58] ), .A(\RF[31][58] ), .S(n10616), .Y(n10276)
         );
  MUX2X1 U13146 ( .B(\RF[28][58] ), .A(\RF[29][58] ), .S(n10616), .Y(n10275)
         );
  MUX2X1 U13147 ( .B(\RF[26][58] ), .A(\RF[27][58] ), .S(n10616), .Y(n10279)
         );
  MUX2X1 U13148 ( .B(\RF[24][58] ), .A(\RF[25][58] ), .S(n10616), .Y(n10278)
         );
  MUX2X1 U13149 ( .B(n10277), .A(n10274), .S(n10693), .Y(n10288) );
  MUX2X1 U13150 ( .B(\RF[22][58] ), .A(\RF[23][58] ), .S(n10616), .Y(n10282)
         );
  MUX2X1 U13151 ( .B(\RF[20][58] ), .A(\RF[21][58] ), .S(n10616), .Y(n10281)
         );
  MUX2X1 U13152 ( .B(\RF[18][58] ), .A(\RF[19][58] ), .S(n10616), .Y(n10285)
         );
  MUX2X1 U13153 ( .B(\RF[16][58] ), .A(\RF[17][58] ), .S(n10616), .Y(n10284)
         );
  MUX2X1 U13154 ( .B(n10283), .A(n10280), .S(n10695), .Y(n10287) );
  MUX2X1 U13155 ( .B(\RF[14][58] ), .A(\RF[15][58] ), .S(n10616), .Y(n10291)
         );
  MUX2X1 U13156 ( .B(\RF[12][58] ), .A(\RF[13][58] ), .S(n10616), .Y(n10290)
         );
  MUX2X1 U13157 ( .B(\RF[10][58] ), .A(\RF[11][58] ), .S(n10616), .Y(n10294)
         );
  MUX2X1 U13158 ( .B(\RF[8][58] ), .A(\RF[9][58] ), .S(n10616), .Y(n10293) );
  MUX2X1 U13159 ( .B(n10292), .A(n10289), .S(n10699), .Y(n10303) );
  MUX2X1 U13160 ( .B(\RF[6][58] ), .A(\RF[7][58] ), .S(n10617), .Y(n10297) );
  MUX2X1 U13161 ( .B(\RF[4][58] ), .A(\RF[5][58] ), .S(n10617), .Y(n10296) );
  MUX2X1 U13162 ( .B(\RF[2][58] ), .A(\RF[3][58] ), .S(n10617), .Y(n10300) );
  MUX2X1 U13163 ( .B(\RF[0][58] ), .A(\RF[1][58] ), .S(n10617), .Y(n10299) );
  MUX2X1 U13164 ( .B(n10298), .A(n10295), .S(n10700), .Y(n10302) );
  MUX2X1 U13165 ( .B(n10301), .A(n10286), .S(N22), .Y(n10512) );
  MUX2X1 U13166 ( .B(\RF[30][59] ), .A(\RF[31][59] ), .S(n10617), .Y(n10306)
         );
  MUX2X1 U13167 ( .B(\RF[28][59] ), .A(\RF[29][59] ), .S(n10617), .Y(n10305)
         );
  MUX2X1 U13168 ( .B(\RF[26][59] ), .A(\RF[27][59] ), .S(n10617), .Y(n10309)
         );
  MUX2X1 U13169 ( .B(\RF[24][59] ), .A(\RF[25][59] ), .S(n10617), .Y(n10308)
         );
  MUX2X1 U13170 ( .B(n10307), .A(n10304), .S(n10684), .Y(n10318) );
  MUX2X1 U13171 ( .B(\RF[22][59] ), .A(\RF[23][59] ), .S(n10617), .Y(n10312)
         );
  MUX2X1 U13172 ( .B(\RF[20][59] ), .A(\RF[21][59] ), .S(n10617), .Y(n10311)
         );
  MUX2X1 U13173 ( .B(\RF[18][59] ), .A(\RF[19][59] ), .S(n10617), .Y(n10315)
         );
  MUX2X1 U13174 ( .B(\RF[16][59] ), .A(\RF[17][59] ), .S(n10617), .Y(n10314)
         );
  MUX2X1 U13175 ( .B(n10313), .A(n10310), .S(n10685), .Y(n10317) );
  MUX2X1 U13176 ( .B(\RF[14][59] ), .A(\RF[15][59] ), .S(n10618), .Y(n10321)
         );
  MUX2X1 U13177 ( .B(\RF[12][59] ), .A(\RF[13][59] ), .S(n10618), .Y(n10320)
         );
  MUX2X1 U13178 ( .B(\RF[10][59] ), .A(\RF[11][59] ), .S(n10618), .Y(n10324)
         );
  MUX2X1 U13179 ( .B(\RF[8][59] ), .A(\RF[9][59] ), .S(n10618), .Y(n10323) );
  MUX2X1 U13180 ( .B(n10322), .A(n10319), .S(n10694), .Y(n10333) );
  MUX2X1 U13181 ( .B(\RF[6][59] ), .A(\RF[7][59] ), .S(n10618), .Y(n10327) );
  MUX2X1 U13182 ( .B(\RF[4][59] ), .A(\RF[5][59] ), .S(n10618), .Y(n10326) );
  MUX2X1 U13183 ( .B(\RF[2][59] ), .A(\RF[3][59] ), .S(n10618), .Y(n10330) );
  MUX2X1 U13184 ( .B(\RF[0][59] ), .A(\RF[1][59] ), .S(n10618), .Y(n10329) );
  MUX2X1 U13185 ( .B(n10328), .A(n10325), .S(n10685), .Y(n10332) );
  MUX2X1 U13186 ( .B(n10331), .A(n10316), .S(N22), .Y(n10513) );
  MUX2X1 U13187 ( .B(\RF[30][60] ), .A(\RF[31][60] ), .S(n10618), .Y(n10336)
         );
  MUX2X1 U13188 ( .B(\RF[28][60] ), .A(\RF[29][60] ), .S(n10618), .Y(n10335)
         );
  MUX2X1 U13189 ( .B(\RF[26][60] ), .A(\RF[27][60] ), .S(n10618), .Y(n10339)
         );
  MUX2X1 U13190 ( .B(\RF[24][60] ), .A(\RF[25][60] ), .S(n10618), .Y(n10338)
         );
  MUX2X1 U13191 ( .B(n10337), .A(n10334), .S(n10688), .Y(n10348) );
  MUX2X1 U13192 ( .B(\RF[22][60] ), .A(\RF[23][60] ), .S(n10619), .Y(n10342)
         );
  MUX2X1 U13193 ( .B(\RF[20][60] ), .A(\RF[21][60] ), .S(n10619), .Y(n10341)
         );
  MUX2X1 U13194 ( .B(\RF[18][60] ), .A(\RF[19][60] ), .S(n10619), .Y(n10345)
         );
  MUX2X1 U13195 ( .B(\RF[16][60] ), .A(\RF[17][60] ), .S(n10619), .Y(n10344)
         );
  MUX2X1 U13196 ( .B(n10343), .A(n10340), .S(n10690), .Y(n10347) );
  MUX2X1 U13197 ( .B(\RF[14][60] ), .A(\RF[15][60] ), .S(n10619), .Y(n10351)
         );
  MUX2X1 U13198 ( .B(\RF[12][60] ), .A(\RF[13][60] ), .S(n10619), .Y(n10350)
         );
  MUX2X1 U13199 ( .B(\RF[10][60] ), .A(\RF[11][60] ), .S(n10619), .Y(n10354)
         );
  MUX2X1 U13200 ( .B(\RF[8][60] ), .A(\RF[9][60] ), .S(n10619), .Y(n10353) );
  MUX2X1 U13201 ( .B(n10352), .A(n10349), .S(n10691), .Y(n10363) );
  MUX2X1 U13202 ( .B(\RF[6][60] ), .A(\RF[7][60] ), .S(n10619), .Y(n10357) );
  MUX2X1 U13203 ( .B(\RF[4][60] ), .A(\RF[5][60] ), .S(n10619), .Y(n10356) );
  MUX2X1 U13204 ( .B(\RF[2][60] ), .A(\RF[3][60] ), .S(n10619), .Y(n10360) );
  MUX2X1 U13205 ( .B(\RF[0][60] ), .A(\RF[1][60] ), .S(n10619), .Y(n10359) );
  MUX2X1 U13206 ( .B(n10358), .A(n10355), .S(n10696), .Y(n10362) );
  MUX2X1 U13207 ( .B(n10361), .A(n10346), .S(N22), .Y(n10514) );
  MUX2X1 U13208 ( .B(\RF[30][61] ), .A(\RF[31][61] ), .S(n10620), .Y(n10366)
         );
  MUX2X1 U13209 ( .B(\RF[28][61] ), .A(\RF[29][61] ), .S(n10620), .Y(n10365)
         );
  MUX2X1 U13210 ( .B(\RF[26][61] ), .A(\RF[27][61] ), .S(n10620), .Y(n10369)
         );
  MUX2X1 U13211 ( .B(\RF[24][61] ), .A(\RF[25][61] ), .S(n10620), .Y(n10368)
         );
  MUX2X1 U13212 ( .B(n10367), .A(n10364), .S(N20), .Y(n10378) );
  MUX2X1 U13213 ( .B(\RF[22][61] ), .A(\RF[23][61] ), .S(n10620), .Y(n10372)
         );
  MUX2X1 U13214 ( .B(\RF[20][61] ), .A(\RF[21][61] ), .S(n10620), .Y(n10371)
         );
  MUX2X1 U13215 ( .B(\RF[18][61] ), .A(\RF[19][61] ), .S(n10620), .Y(n10375)
         );
  MUX2X1 U13216 ( .B(\RF[16][61] ), .A(\RF[17][61] ), .S(n10620), .Y(n10374)
         );
  MUX2X1 U13217 ( .B(n10373), .A(n10370), .S(N20), .Y(n10377) );
  MUX2X1 U13218 ( .B(\RF[14][61] ), .A(\RF[15][61] ), .S(n10620), .Y(n10381)
         );
  MUX2X1 U13219 ( .B(\RF[12][61] ), .A(\RF[13][61] ), .S(n10620), .Y(n10380)
         );
  MUX2X1 U13220 ( .B(\RF[10][61] ), .A(\RF[11][61] ), .S(n10620), .Y(n10384)
         );
  MUX2X1 U13221 ( .B(\RF[8][61] ), .A(\RF[9][61] ), .S(n10620), .Y(n10383) );
  MUX2X1 U13222 ( .B(n10382), .A(n10379), .S(N20), .Y(n10393) );
  MUX2X1 U13223 ( .B(\RF[6][61] ), .A(\RF[7][61] ), .S(n10621), .Y(n10387) );
  MUX2X1 U13224 ( .B(\RF[4][61] ), .A(\RF[5][61] ), .S(n10621), .Y(n10386) );
  MUX2X1 U13225 ( .B(\RF[2][61] ), .A(\RF[3][61] ), .S(n10621), .Y(n10390) );
  MUX2X1 U13226 ( .B(\RF[0][61] ), .A(\RF[1][61] ), .S(n10621), .Y(n10389) );
  MUX2X1 U13227 ( .B(n10388), .A(n10385), .S(N20), .Y(n10392) );
  MUX2X1 U13228 ( .B(n10391), .A(n10376), .S(N22), .Y(n10515) );
  MUX2X1 U13229 ( .B(\RF[30][62] ), .A(\RF[31][62] ), .S(n10621), .Y(n10396)
         );
  MUX2X1 U13230 ( .B(\RF[28][62] ), .A(\RF[29][62] ), .S(n10621), .Y(n10395)
         );
  MUX2X1 U13231 ( .B(\RF[26][62] ), .A(\RF[27][62] ), .S(n10621), .Y(n10399)
         );
  MUX2X1 U13232 ( .B(\RF[24][62] ), .A(\RF[25][62] ), .S(n10621), .Y(n10398)
         );
  MUX2X1 U13233 ( .B(n10397), .A(n10394), .S(N20), .Y(n10408) );
  MUX2X1 U13234 ( .B(\RF[22][62] ), .A(\RF[23][62] ), .S(n10621), .Y(n10402)
         );
  MUX2X1 U13235 ( .B(\RF[20][62] ), .A(\RF[21][62] ), .S(n10621), .Y(n10401)
         );
  MUX2X1 U13236 ( .B(\RF[18][62] ), .A(\RF[19][62] ), .S(n10621), .Y(n10405)
         );
  MUX2X1 U13237 ( .B(\RF[16][62] ), .A(\RF[17][62] ), .S(n10621), .Y(n10404)
         );
  MUX2X1 U13238 ( .B(n10403), .A(n10400), .S(N20), .Y(n10407) );
  MUX2X1 U13239 ( .B(\RF[14][62] ), .A(\RF[15][62] ), .S(n10622), .Y(n10411)
         );
  MUX2X1 U13240 ( .B(\RF[12][62] ), .A(\RF[13][62] ), .S(n10622), .Y(n10410)
         );
  MUX2X1 U13241 ( .B(\RF[10][62] ), .A(\RF[11][62] ), .S(n10622), .Y(n10414)
         );
  MUX2X1 U13242 ( .B(\RF[8][62] ), .A(\RF[9][62] ), .S(n10622), .Y(n10413) );
  MUX2X1 U13243 ( .B(n10412), .A(n10409), .S(N20), .Y(n10423) );
  MUX2X1 U13244 ( .B(\RF[6][62] ), .A(\RF[7][62] ), .S(n10622), .Y(n10417) );
  MUX2X1 U13245 ( .B(\RF[4][62] ), .A(\RF[5][62] ), .S(n10622), .Y(n10416) );
  MUX2X1 U13246 ( .B(\RF[2][62] ), .A(\RF[3][62] ), .S(n10622), .Y(n10420) );
  MUX2X1 U13247 ( .B(\RF[0][62] ), .A(\RF[1][62] ), .S(n10622), .Y(n10419) );
  MUX2X1 U13248 ( .B(n10418), .A(n10415), .S(N20), .Y(n10422) );
  MUX2X1 U13249 ( .B(n10421), .A(n10406), .S(N22), .Y(n10516) );
  MUX2X1 U13250 ( .B(\RF[30][63] ), .A(\RF[31][63] ), .S(n10622), .Y(n10426)
         );
  MUX2X1 U13251 ( .B(\RF[28][63] ), .A(\RF[29][63] ), .S(n10622), .Y(n10425)
         );
  MUX2X1 U13252 ( .B(\RF[26][63] ), .A(\RF[27][63] ), .S(n10622), .Y(n10429)
         );
  MUX2X1 U13253 ( .B(\RF[24][63] ), .A(\RF[25][63] ), .S(n10622), .Y(n10428)
         );
  MUX2X1 U13254 ( .B(n10427), .A(n10424), .S(n10692), .Y(n10438) );
  MUX2X1 U13255 ( .B(\RF[22][63] ), .A(\RF[23][63] ), .S(n10623), .Y(n10432)
         );
  MUX2X1 U13256 ( .B(\RF[20][63] ), .A(\RF[21][63] ), .S(n10623), .Y(n10431)
         );
  MUX2X1 U13257 ( .B(\RF[18][63] ), .A(\RF[19][63] ), .S(n10623), .Y(n10435)
         );
  MUX2X1 U13258 ( .B(\RF[16][63] ), .A(\RF[17][63] ), .S(n10623), .Y(n10434)
         );
  MUX2X1 U13259 ( .B(n10433), .A(n10430), .S(n10697), .Y(n10437) );
  MUX2X1 U13260 ( .B(\RF[14][63] ), .A(\RF[15][63] ), .S(n10623), .Y(n10441)
         );
  MUX2X1 U13261 ( .B(\RF[12][63] ), .A(\RF[13][63] ), .S(n10623), .Y(n10440)
         );
  MUX2X1 U13262 ( .B(\RF[10][63] ), .A(\RF[11][63] ), .S(n10623), .Y(n10444)
         );
  MUX2X1 U13263 ( .B(\RF[8][63] ), .A(\RF[9][63] ), .S(n10623), .Y(n10443) );
  MUX2X1 U13264 ( .B(n10442), .A(n10439), .S(n10689), .Y(n10453) );
  MUX2X1 U13265 ( .B(\RF[6][63] ), .A(\RF[7][63] ), .S(n10623), .Y(n10447) );
  MUX2X1 U13266 ( .B(\RF[4][63] ), .A(\RF[5][63] ), .S(n10623), .Y(n10446) );
  MUX2X1 U13267 ( .B(\RF[2][63] ), .A(\RF[3][63] ), .S(n10623), .Y(n10450) );
  MUX2X1 U13268 ( .B(\RF[0][63] ), .A(\RF[1][63] ), .S(n10623), .Y(n10449) );
  MUX2X1 U13269 ( .B(n10448), .A(n10445), .S(n10698), .Y(n10452) );
  MUX2X1 U13270 ( .B(n10451), .A(n10436), .S(N22), .Y(n10517) );
endmodule

